module tt_um_dlfloatmac (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \MAC.a[0] ;
 wire \MAC.a[10] ;
 wire \MAC.a[11] ;
 wire \MAC.a[12] ;
 wire \MAC.a[13] ;
 wire \MAC.a[14] ;
 wire \MAC.a[15] ;
 wire \MAC.a[1] ;
 wire \MAC.a[2] ;
 wire \MAC.a[3] ;
 wire \MAC.a[4] ;
 wire \MAC.a[5] ;
 wire \MAC.a[6] ;
 wire \MAC.a[7] ;
 wire \MAC.a[8] ;
 wire \MAC.a[9] ;
 wire \MAC.add.a1[0] ;
 wire \MAC.add.a1[10] ;
 wire \MAC.add.a1[11] ;
 wire \MAC.add.a1[12] ;
 wire \MAC.add.a1[13] ;
 wire \MAC.add.a1[14] ;
 wire \MAC.add.a1[15] ;
 wire \MAC.add.a1[1] ;
 wire \MAC.add.a1[2] ;
 wire \MAC.add.a1[3] ;
 wire \MAC.add.a1[4] ;
 wire \MAC.add.a1[5] ;
 wire \MAC.add.a1[6] ;
 wire \MAC.add.a1[7] ;
 wire \MAC.add.a1[8] ;
 wire \MAC.add.a1[9] ;
 wire \MAC.add.b1[0] ;
 wire \MAC.add.b1[10] ;
 wire \MAC.add.b1[11] ;
 wire \MAC.add.b1[12] ;
 wire \MAC.add.b1[13] ;
 wire \MAC.add.b1[14] ;
 wire \MAC.add.b1[15] ;
 wire \MAC.add.b1[1] ;
 wire \MAC.add.b1[2] ;
 wire \MAC.add.b1[3] ;
 wire \MAC.add.b1[4] ;
 wire \MAC.add.b1[5] ;
 wire \MAC.add.b1[6] ;
 wire \MAC.add.b1[7] ;
 wire \MAC.add.b1[8] ;
 wire \MAC.add.b1[9] ;
 wire \MAC.add.c_add[0] ;
 wire \MAC.add.c_add[10] ;
 wire \MAC.add.c_add[11] ;
 wire \MAC.add.c_add[12] ;
 wire \MAC.add.c_add[13] ;
 wire \MAC.add.c_add[14] ;
 wire \MAC.add.c_add[1] ;
 wire \MAC.add.c_add[2] ;
 wire \MAC.add.c_add[3] ;
 wire \MAC.add.c_add[4] ;
 wire \MAC.add.c_add[5] ;
 wire \MAC.add.c_add[6] ;
 wire \MAC.add.c_add[7] ;
 wire \MAC.add.c_add[8] ;
 wire \MAC.add.c_add[9] ;
 wire \MAC.b[0] ;
 wire \MAC.b[10] ;
 wire \MAC.b[11] ;
 wire \MAC.b[12] ;
 wire \MAC.b[13] ;
 wire \MAC.b[14] ;
 wire \MAC.b[15] ;
 wire \MAC.b[1] ;
 wire \MAC.b[2] ;
 wire \MAC.b[3] ;
 wire \MAC.b[4] ;
 wire \MAC.b[5] ;
 wire \MAC.b[6] ;
 wire \MAC.b[7] ;
 wire \MAC.b[8] ;
 wire \MAC.b[9] ;
 wire \MAC.mul.c_mul1[0] ;
 wire \MAC.mul.c_mul1[10] ;
 wire \MAC.mul.c_mul1[11] ;
 wire \MAC.mul.c_mul1[12] ;
 wire \MAC.mul.c_mul1[13] ;
 wire \MAC.mul.c_mul1[14] ;
 wire \MAC.mul.c_mul1[15] ;
 wire \MAC.mul.c_mul1[1] ;
 wire \MAC.mul.c_mul1[2] ;
 wire \MAC.mul.c_mul1[3] ;
 wire \MAC.mul.c_mul1[4] ;
 wire \MAC.mul.c_mul1[5] ;
 wire \MAC.mul.c_mul1[6] ;
 wire \MAC.mul.c_mul1[7] ;
 wire \MAC.mul.c_mul1[8] ;
 wire \MAC.mul.c_mul1[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire clknet_0_clk;
 wire \wrap.state[0] ;
 wire \wrap.temp_data[0] ;
 wire \wrap.temp_data[10] ;
 wire \wrap.temp_data[11] ;
 wire \wrap.temp_data[12] ;
 wire \wrap.temp_data[13] ;
 wire \wrap.temp_data[14] ;
 wire \wrap.temp_data[15] ;
 wire \wrap.temp_data[1] ;
 wire \wrap.temp_data[2] ;
 wire \wrap.temp_data[3] ;
 wire \wrap.temp_data[4] ;
 wire \wrap.temp_data[5] ;
 wire \wrap.temp_data[6] ;
 wire \wrap.temp_data[7] ;
 wire \wrap.temp_data[8] ;
 wire \wrap.temp_data[9] ;
 wire \wrap2.state[0] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;

 sky130_fd_sc_hd__inv_2 _1177_ (.A(\wrap.state[0] ),
    .Y(_0415_));
 sky130_fd_sc_hd__buf_2 _1178_ (.A(_0415_),
    .X(_0000_));
 sky130_fd_sc_hd__inv_2 _1179_ (.A(net47),
    .Y(_0001_));
 sky130_fd_sc_hd__clkbuf_2 _1180_ (.A(\wrap.state[0] ),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _1181_ (.A(_0416_),
    .B(net46),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _1182_ (.A(_0417_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _1183_ (.A(_0416_),
    .B(net54),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _1184_ (.A(_0418_),
    .X(_0009_));
 sky130_fd_sc_hd__and2_1 _1185_ (.A(_0416_),
    .B(net50),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _1186_ (.A(_0419_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_2 _1187_ (.A(\wrap.state[0] ),
    .X(_0420_));
 sky130_fd_sc_hd__and2_1 _1188_ (.A(_0420_),
    .B(net61),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _1189_ (.A(_0421_),
    .X(_0011_));
 sky130_fd_sc_hd__and2_1 _1190_ (.A(_0420_),
    .B(net60),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _1191_ (.A(_0422_),
    .X(_0012_));
 sky130_fd_sc_hd__and2_1 _1192_ (.A(_0420_),
    .B(net56),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _1193_ (.A(_0423_),
    .X(_0013_));
 sky130_fd_sc_hd__and2_1 _1194_ (.A(_0420_),
    .B(net53),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _1195_ (.A(_0424_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _1196_ (.A(_0420_),
    .B(net55),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_1 _1197_ (.A(_0425_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _1198_ (.A(_0420_),
    .B(net52),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_1 _1199_ (.A(_0426_),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _1200_ (.A(_0420_),
    .B(net51),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _1201_ (.A(_0427_),
    .X(_0017_));
 sky130_fd_sc_hd__and2_1 _1202_ (.A(_0420_),
    .B(net48),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_1 _1203_ (.A(_0428_),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _1204_ (.A(_0420_),
    .B(net57),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_1 _1205_ (.A(_0429_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _1206_ (.A(_0420_),
    .B(net58),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _1207_ (.A(_0430_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _1208_ (.A(\wrap.state[0] ),
    .B(net59),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _1209_ (.A(_0431_),
    .X(_0006_));
 sky130_fd_sc_hd__and2_1 _1210_ (.A(\wrap.state[0] ),
    .B(net62),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _1211_ (.A(_0432_),
    .X(_0007_));
 sky130_fd_sc_hd__and2_1 _1212_ (.A(\wrap.state[0] ),
    .B(net49),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _1213_ (.A(_0433_),
    .X(_0008_));
 sky130_fd_sc_hd__clkbuf_2 _1214_ (.A(_0416_),
    .X(_0434_));
 sky130_fd_sc_hd__and2_1 _1215_ (.A(_0434_),
    .B(net2),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _1216_ (.A(_0435_),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _1217_ (.A(_0434_),
    .B(net3),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _1218_ (.A(_0436_),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _1219_ (.A(_0434_),
    .B(net4),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _1220_ (.A(_0437_),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _1221_ (.A(_0434_),
    .B(net5),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _1222_ (.A(_0438_),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _1223_ (.A(_0434_),
    .B(net6),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_1 _1224_ (.A(_0439_),
    .X(_0028_));
 sky130_fd_sc_hd__and2_1 _1225_ (.A(_0434_),
    .B(net7),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_1 _1226_ (.A(_0440_),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _1227_ (.A(_0434_),
    .B(net8),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_1 _1228_ (.A(_0441_),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _1229_ (.A(_0434_),
    .B(net9),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _1230_ (.A(_0442_),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _1231_ (.A(_0434_),
    .B(net10),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _1232_ (.A(_0443_),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _1233_ (.A(_0434_),
    .B(net11),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _1234_ (.A(_0444_),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _1235_ (.A(_0416_),
    .B(net12),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _1236_ (.A(_0445_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _1237_ (.A(_0416_),
    .B(net13),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _1238_ (.A(_0446_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _1239_ (.A(_0416_),
    .B(net14),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _1240_ (.A(_0447_),
    .X(_0021_));
 sky130_fd_sc_hd__and2_1 _1241_ (.A(_0416_),
    .B(net15),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _1242_ (.A(_0448_),
    .X(_0022_));
 sky130_fd_sc_hd__and2_1 _1243_ (.A(_0416_),
    .B(net16),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _1244_ (.A(_0449_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _1245_ (.A(_0416_),
    .B(net17),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _1246_ (.A(_0450_),
    .X(_0024_));
 sky130_fd_sc_hd__or4_1 _1247_ (.A(\MAC.add.a1[12] ),
    .B(\MAC.add.a1[11] ),
    .C(\MAC.add.a1[10] ),
    .D(\MAC.add.a1[9] ),
    .X(_0451_));
 sky130_fd_sc_hd__nor3_1 _1248_ (.A(\MAC.add.a1[14] ),
    .B(\MAC.add.a1[13] ),
    .C(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__or4_1 _1249_ (.A(\MAC.add.b1[12] ),
    .B(\MAC.add.b1[11] ),
    .C(\MAC.add.b1[10] ),
    .D(\MAC.add.b1[9] ),
    .X(_0453_));
 sky130_fd_sc_hd__nor3_1 _1250_ (.A(\MAC.add.b1[14] ),
    .B(\MAC.add.b1[13] ),
    .C(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__or2_1 _1251_ (.A(_0452_),
    .B(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_4 _1252_ (.A(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__buf_2 _1253_ (.A(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__or2b_2 _1254_ (.A(\MAC.add.a1[14] ),
    .B_N(\MAC.add.b1[14] ),
    .X(_0458_));
 sky130_fd_sc_hd__and2b_1 _1255_ (.A_N(\MAC.add.b1[13] ),
    .B(\MAC.add.a1[13] ),
    .X(_0459_));
 sky130_fd_sc_hd__and2b_1 _1256_ (.A_N(\MAC.add.a1[13] ),
    .B(\MAC.add.b1[13] ),
    .X(_0460_));
 sky130_fd_sc_hd__nor2_1 _1257_ (.A(_0459_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__inv_2 _1258_ (.A(\MAC.add.b1[12] ),
    .Y(_0462_));
 sky130_fd_sc_hd__xnor2_2 _1259_ (.A(\MAC.add.b1[10] ),
    .B(\MAC.add.a1[10] ),
    .Y(_0463_));
 sky130_fd_sc_hd__or2b_1 _1260_ (.A(\MAC.add.a1[9] ),
    .B_N(\MAC.add.b1[9] ),
    .X(_0464_));
 sky130_fd_sc_hd__and2b_1 _1261_ (.A_N(\MAC.add.b1[10] ),
    .B(\MAC.add.a1[10] ),
    .X(_0465_));
 sky130_fd_sc_hd__a21o_1 _1262_ (.A1(_0463_),
    .A2(_0464_),
    .B1(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__xnor2_2 _1263_ (.A(\MAC.add.b1[12] ),
    .B(\MAC.add.a1[12] ),
    .Y(_0467_));
 sky130_fd_sc_hd__xnor2_2 _1264_ (.A(\MAC.add.b1[11] ),
    .B(\MAC.add.a1[11] ),
    .Y(_0468_));
 sky130_fd_sc_hd__and2_1 _1265_ (.A(_0467_),
    .B(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__and2b_1 _1266_ (.A_N(\MAC.add.b1[11] ),
    .B(\MAC.add.a1[11] ),
    .X(_0470_));
 sky130_fd_sc_hd__o21a_1 _1267_ (.A1(_0462_),
    .A2(\MAC.add.a1[12] ),
    .B1(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__a221o_1 _1268_ (.A1(_0462_),
    .A2(\MAC.add.a1[12] ),
    .B1(_0466_),
    .B2(_0469_),
    .C1(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__and2b_1 _1269_ (.A_N(\MAC.add.b1[14] ),
    .B(\MAC.add.a1[14] ),
    .X(_0473_));
 sky130_fd_sc_hd__a211o_4 _1270_ (.A1(_0472_),
    .A2(_0461_),
    .B1(_0473_),
    .C1(_0459_),
    .X(_0474_));
 sky130_fd_sc_hd__xnor2_2 _1271_ (.A(\MAC.add.b1[9] ),
    .B(\MAC.add.a1[9] ),
    .Y(_0475_));
 sky130_fd_sc_hd__and2_1 _1272_ (.A(_0463_),
    .B(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__nand3_1 _1273_ (.A(_0467_),
    .B(_0468_),
    .C(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__or3b_4 _1274_ (.A(_0477_),
    .B(_0473_),
    .C_N(_0461_),
    .X(_0478_));
 sky130_fd_sc_hd__nand3_4 _1275_ (.A(_0458_),
    .B(_0474_),
    .C(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__a21oi_1 _1276_ (.A1(_0466_),
    .A2(_0468_),
    .B1(_0470_),
    .Y(_0480_));
 sky130_fd_sc_hd__xnor2_1 _1277_ (.A(_0467_),
    .B(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__buf_2 _1278_ (.A(_0458_),
    .X(_0482_));
 sky130_fd_sc_hd__buf_2 _1279_ (.A(_0474_),
    .X(_0483_));
 sky130_fd_sc_hd__buf_2 _1280_ (.A(_0478_),
    .X(_0484_));
 sky130_fd_sc_hd__or2b_1 _1281_ (.A(\MAC.add.a1[11] ),
    .B_N(\MAC.add.b1[11] ),
    .X(_0485_));
 sky130_fd_sc_hd__nand2_1 _1282_ (.A(_0463_),
    .B(_0475_),
    .Y(_0486_));
 sky130_fd_sc_hd__a31o_1 _1283_ (.A1(_0466_),
    .A2(_0485_),
    .A3(_0486_),
    .B1(_0470_),
    .X(_0487_));
 sky130_fd_sc_hd__xnor2_1 _1284_ (.A(_0467_),
    .B(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__a31o_1 _1285_ (.A1(_0482_),
    .A2(_0483_),
    .A3(_0484_),
    .B1(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nor2_1 _1286_ (.A(_0452_),
    .B(_0454_),
    .Y(_0490_));
 sky130_fd_sc_hd__clkbuf_4 _1287_ (.A(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__o211a_1 _1288_ (.A1(_0479_),
    .A2(_0481_),
    .B1(_0489_),
    .C1(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__xor2_1 _1289_ (.A(_0461_),
    .B(_0472_),
    .X(_0493_));
 sky130_fd_sc_hd__and2b_1 _1290_ (.A_N(\MAC.add.a1[14] ),
    .B(\MAC.add.b1[14] ),
    .X(_0494_));
 sky130_fd_sc_hd__a21oi_1 _1291_ (.A1(_0461_),
    .A2(_0472_),
    .B1(_0459_),
    .Y(_0495_));
 sky130_fd_sc_hd__or2b_1 _1292_ (.A(\MAC.add.b1[14] ),
    .B_N(\MAC.add.a1[14] ),
    .X(_0496_));
 sky130_fd_sc_hd__o211a_1 _1293_ (.A1(_0494_),
    .A2(_0495_),
    .B1(_0477_),
    .C1(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__o2111ai_1 _1294_ (.A1(_0494_),
    .A2(_0495_),
    .B1(_0477_),
    .C1(_0493_),
    .D1(_0496_),
    .Y(_0498_));
 sky130_fd_sc_hd__o211a_1 _1295_ (.A1(_0493_),
    .A2(_0497_),
    .B1(_0498_),
    .C1(_0491_),
    .X(_0499_));
 sky130_fd_sc_hd__nor2_1 _1296_ (.A(_0492_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__xnor2_1 _1297_ (.A(_0463_),
    .B(_0464_),
    .Y(_0501_));
 sky130_fd_sc_hd__a31o_1 _1298_ (.A1(_0482_),
    .A2(_0483_),
    .A3(_0484_),
    .B1(_0475_),
    .X(_0502_));
 sky130_fd_sc_hd__a311oi_1 _1299_ (.A1(_0482_),
    .A2(_0483_),
    .A3(_0484_),
    .B1(_0501_),
    .C1(_0475_),
    .Y(_0503_));
 sky130_fd_sc_hd__a211oi_2 _1300_ (.A1(_0501_),
    .A2(_0502_),
    .B1(_0503_),
    .C1(_0456_),
    .Y(_0504_));
 sky130_fd_sc_hd__o21ai_2 _1301_ (.A1(_0494_),
    .A2(_0478_),
    .B1(_0490_),
    .Y(_0505_));
 sky130_fd_sc_hd__clkbuf_4 _1302_ (.A(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__a211o_1 _1303_ (.A1(_0461_),
    .A2(_0472_),
    .B1(_0458_),
    .C1(_0459_),
    .X(_0507_));
 sky130_fd_sc_hd__o211a_2 _1304_ (.A1(_0496_),
    .A2(_0495_),
    .B1(_0478_),
    .C1(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__or2_1 _1305_ (.A(_0506_),
    .B(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__nor2_2 _1306_ (.A(_0475_),
    .B(_0456_),
    .Y(_0510_));
 sky130_fd_sc_hd__a31o_1 _1307_ (.A1(_0482_),
    .A2(_0483_),
    .A3(_0484_),
    .B1(\MAC.add.a1[8] ),
    .X(_0511_));
 sky130_fd_sc_hd__o221a_1 _1308_ (.A1(\MAC.add.b1[8] ),
    .A2(_0479_),
    .B1(_0506_),
    .B2(_0508_),
    .C1(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__a21oi_1 _1309_ (.A1(_0509_),
    .A2(_0510_),
    .B1(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__or2_1 _1310_ (.A(net18),
    .B(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__xnor2_1 _1311_ (.A(_0466_),
    .B(_0468_),
    .Y(_0515_));
 sky130_fd_sc_hd__a31o_1 _1312_ (.A1(_0458_),
    .A2(_0474_),
    .A3(_0484_),
    .B1(_0476_),
    .X(_0516_));
 sky130_fd_sc_hd__xnor2_1 _1313_ (.A(_0515_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__nor2_1 _1314_ (.A(_0456_),
    .B(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__nor2_1 _1315_ (.A(_0499_),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__and2b_1 _1316_ (.A_N(_0514_),
    .B(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__or2_1 _1317_ (.A(_0456_),
    .B(_0517_),
    .X(_0521_));
 sky130_fd_sc_hd__a31o_1 _1318_ (.A1(_0482_),
    .A2(_0483_),
    .A3(_0484_),
    .B1(\MAC.add.a1[5] ),
    .X(_0522_));
 sky130_fd_sc_hd__o221a_1 _1319_ (.A1(\MAC.add.b1[5] ),
    .A2(_0479_),
    .B1(_0505_),
    .B2(_0508_),
    .C1(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__a31o_1 _1320_ (.A1(_0482_),
    .A2(_0483_),
    .A3(_0484_),
    .B1(\MAC.add.a1[4] ),
    .X(_0524_));
 sky130_fd_sc_hd__o221a_1 _1321_ (.A1(\MAC.add.b1[4] ),
    .A2(_0479_),
    .B1(_0505_),
    .B2(_0508_),
    .C1(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__or2_2 _1322_ (.A(_0475_),
    .B(_0455_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _1323_ (.A0(_0523_),
    .A1(_0525_),
    .S(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__a31o_1 _1324_ (.A1(_0482_),
    .A2(_0483_),
    .A3(_0484_),
    .B1(\MAC.add.a1[7] ),
    .X(_0528_));
 sky130_fd_sc_hd__o221a_1 _1325_ (.A1(\MAC.add.b1[7] ),
    .A2(_0479_),
    .B1(_0505_),
    .B2(_0508_),
    .C1(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__a31o_1 _1326_ (.A1(_0482_),
    .A2(_0483_),
    .A3(_0484_),
    .B1(\MAC.add.a1[6] ),
    .X(_0530_));
 sky130_fd_sc_hd__o221a_1 _1327_ (.A1(\MAC.add.b1[6] ),
    .A2(_0479_),
    .B1(_0505_),
    .B2(_0508_),
    .C1(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _1328_ (.A0(_0529_),
    .A1(_0531_),
    .S(_0526_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _1329_ (.A0(_0527_),
    .A1(_0532_),
    .S(net18),
    .X(_0533_));
 sky130_fd_sc_hd__a211o_1 _1330_ (.A1(_0501_),
    .A2(_0502_),
    .B1(_0503_),
    .C1(_0455_),
    .X(_0534_));
 sky130_fd_sc_hd__o21a_1 _1331_ (.A1(_0506_),
    .A2(_0508_),
    .B1(_0526_),
    .X(_0535_));
 sky130_fd_sc_hd__and2_1 _1332_ (.A(_0534_),
    .B(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__and3_1 _1333_ (.A(_0458_),
    .B(_0474_),
    .C(_0478_),
    .X(_0537_));
 sky130_fd_sc_hd__clkbuf_4 _1334_ (.A(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _1335_ (.A0(\MAC.add.a1[0] ),
    .A1(\MAC.add.b1[0] ),
    .S(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__a21o_1 _1336_ (.A1(_0536_),
    .A2(_0539_),
    .B1(_0518_),
    .X(_0540_));
 sky130_fd_sc_hd__a31o_1 _1337_ (.A1(_0482_),
    .A2(_0483_),
    .A3(_0484_),
    .B1(\MAC.add.a1[3] ),
    .X(_0541_));
 sky130_fd_sc_hd__o221a_1 _1338_ (.A1(\MAC.add.b1[3] ),
    .A2(_0479_),
    .B1(_0506_),
    .B2(_0508_),
    .C1(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _1339_ (.A0(\MAC.add.a1[2] ),
    .A1(\MAC.add.b1[2] ),
    .S(_0538_),
    .X(_0543_));
 sky130_fd_sc_hd__a22o_1 _1340_ (.A1(_0510_),
    .A2(_0542_),
    .B1(_0543_),
    .B2(_0535_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _1341_ (.A0(\MAC.add.a1[1] ),
    .A1(\MAC.add.b1[1] ),
    .S(_0538_),
    .X(_0545_));
 sky130_fd_sc_hd__and3_1 _1342_ (.A(_0509_),
    .B(_0510_),
    .C(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _1343_ (.A0(_0544_),
    .A1(_0546_),
    .S(_0534_),
    .X(_0547_));
 sky130_fd_sc_hd__o22a_1 _1344_ (.A1(_0521_),
    .A2(_0533_),
    .B1(_0540_),
    .B2(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__o22a_1 _1345_ (.A1(_0500_),
    .A2(_0520_),
    .B1(_0548_),
    .B2(_0492_),
    .X(_0549_));
 sky130_fd_sc_hd__inv_2 _1346_ (.A(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__inv_2 _1347_ (.A(\MAC.add.a1[0] ),
    .Y(_0551_));
 sky130_fd_sc_hd__inv_2 _1348_ (.A(\MAC.add.b1[0] ),
    .Y(_0552_));
 sky130_fd_sc_hd__clkbuf_4 _1349_ (.A(_0479_),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _1350_ (.A0(_0551_),
    .A1(_0552_),
    .S(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__nor2_1 _1351_ (.A(_0550_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__and4_1 _1352_ (.A(_0534_),
    .B(_0509_),
    .C(_0510_),
    .D(_0543_),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _1353_ (.A0(_0542_),
    .A1(_0525_),
    .S(_0510_),
    .X(_0557_));
 sky130_fd_sc_hd__a22o_1 _1354_ (.A1(_0536_),
    .A2(_0545_),
    .B1(_0557_),
    .B2(_0504_),
    .X(_0558_));
 sky130_fd_sc_hd__o21ai_1 _1355_ (.A1(_0556_),
    .A2(_0558_),
    .B1(_0521_),
    .Y(_0559_));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(_0523_),
    .A1(_0531_),
    .S(_0510_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _1357_ (.A0(_0512_),
    .A1(_0529_),
    .S(_0526_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _1358_ (.A0(_0560_),
    .A1(_0561_),
    .S(net18),
    .X(_0562_));
 sky130_fd_sc_hd__a21oi_1 _1359_ (.A1(_0518_),
    .A2(_0562_),
    .B1(_0492_),
    .Y(_0563_));
 sky130_fd_sc_hd__a21oi_1 _1360_ (.A1(_0519_),
    .A2(_0536_),
    .B1(_0500_),
    .Y(_0564_));
 sky130_fd_sc_hd__a21oi_2 _1361_ (.A1(_0559_),
    .A2(_0563_),
    .B1(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__mux2_1 _1362_ (.A0(\MAC.add.a1[1] ),
    .A1(\MAC.add.b1[1] ),
    .S(_0553_),
    .X(_0566_));
 sky130_fd_sc_hd__xnor2_2 _1363_ (.A(\MAC.add.b1[8] ),
    .B(\MAC.add.a1[8] ),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _1364_ (.A(_0534_),
    .B(_0532_),
    .Y(_0568_));
 sky130_fd_sc_hd__o21a_1 _1365_ (.A1(_0534_),
    .A2(_0513_),
    .B1(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__nand2_1 _1366_ (.A(_0500_),
    .B(_0518_),
    .Y(_0570_));
 sky130_fd_sc_hd__and2_1 _1367_ (.A(_0500_),
    .B(_0521_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _1368_ (.A0(_0544_),
    .A1(_0527_),
    .S(net18),
    .X(_0572_));
 sky130_fd_sc_hd__a2bb2o_1 _1369_ (.A1_N(_0569_),
    .A2_N(_0570_),
    .B1(_0571_),
    .B2(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _1370_ (.A0(\MAC.add.a1[2] ),
    .A1(\MAC.add.b1[2] ),
    .S(_0553_),
    .X(_0574_));
 sky130_fd_sc_hd__inv_2 _1371_ (.A(_0574_),
    .Y(_0575_));
 sky130_fd_sc_hd__inv_2 _1372_ (.A(\MAC.add.a1[1] ),
    .Y(_0576_));
 sky130_fd_sc_hd__inv_2 _1373_ (.A(\MAC.add.b1[1] ),
    .Y(_0577_));
 sky130_fd_sc_hd__mux2_1 _1374_ (.A0(_0576_),
    .A1(_0577_),
    .S(_0553_),
    .X(_0578_));
 sky130_fd_sc_hd__o22a_1 _1375_ (.A1(_0565_),
    .A2(_0578_),
    .B1(_0573_),
    .B2(_0575_),
    .X(_0579_));
 sky130_fd_sc_hd__a211o_1 _1376_ (.A1(_0565_),
    .A2(_0578_),
    .B1(_0554_),
    .C1(_0549_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _1377_ (.A0(_0557_),
    .A1(_0560_),
    .S(net18),
    .X(_0581_));
 sky130_fd_sc_hd__nand2_1 _1378_ (.A(_0509_),
    .B(_0526_),
    .Y(_0582_));
 sky130_fd_sc_hd__nor2_1 _1379_ (.A(net18),
    .B(_0561_),
    .Y(_0583_));
 sky130_fd_sc_hd__a21o_1 _1380_ (.A1(net18),
    .A2(_0582_),
    .B1(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__o2bb2a_1 _1381_ (.A1_N(_0581_),
    .A2_N(_0571_),
    .B1(_0570_),
    .B2(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _1382_ (.A0(\MAC.add.a1[3] ),
    .A1(\MAC.add.b1[3] ),
    .S(_0553_),
    .X(_0586_));
 sky130_fd_sc_hd__nor2_1 _1383_ (.A(_0585_),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__a221o_1 _1384_ (.A1(_0573_),
    .A2(_0575_),
    .B1(_0579_),
    .B2(_0580_),
    .C1(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _1385_ (.A0(\MAC.add.a1[5] ),
    .A1(\MAC.add.b1[5] ),
    .S(_0553_),
    .X(_0589_));
 sky130_fd_sc_hd__inv_2 _1386_ (.A(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__and3_1 _1387_ (.A(_0500_),
    .B(_0518_),
    .C(_0536_),
    .X(_0591_));
 sky130_fd_sc_hd__a21o_1 _1388_ (.A1(_0562_),
    .A2(_0571_),
    .B1(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _1389_ (.A0(\MAC.add.a1[4] ),
    .A1(\MAC.add.b1[4] ),
    .S(_0553_),
    .X(_0593_));
 sky130_fd_sc_hd__o2bb2a_1 _1390_ (.A1_N(_0533_),
    .A2_N(_0571_),
    .B1(_0570_),
    .B2(_0514_),
    .X(_0594_));
 sky130_fd_sc_hd__o2bb2a_1 _1391_ (.A1_N(_0590_),
    .A2_N(_0592_),
    .B1(_0593_),
    .B2(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__nand2_1 _1392_ (.A(_0500_),
    .B(_0521_),
    .Y(_0596_));
 sky130_fd_sc_hd__nor2_1 _1393_ (.A(_0596_),
    .B(_0584_),
    .Y(_0597_));
 sky130_fd_sc_hd__mux2_2 _1394_ (.A0(\MAC.add.a1[7] ),
    .A1(\MAC.add.b1[7] ),
    .S(_0553_),
    .X(_0598_));
 sky130_fd_sc_hd__inv_2 _1395_ (.A(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__nor2_1 _1396_ (.A(_0569_),
    .B(_0596_),
    .Y(_0600_));
 sky130_fd_sc_hd__mux2_2 _1397_ (.A0(\MAC.add.a1[6] ),
    .A1(\MAC.add.b1[6] ),
    .S(_0553_),
    .X(_0601_));
 sky130_fd_sc_hd__inv_2 _1398_ (.A(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__a211o_1 _1399_ (.A1(net18),
    .A2(_0582_),
    .B1(_0596_),
    .C1(_0583_),
    .X(_0603_));
 sky130_fd_sc_hd__o32a_1 _1400_ (.A1(_0569_),
    .A2(_0596_),
    .A3(_0601_),
    .B1(_0598_),
    .B2(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__o221a_1 _1401_ (.A1(_0597_),
    .A2(_0599_),
    .B1(_0600_),
    .B2(_0602_),
    .C1(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__or2_1 _1402_ (.A(_0592_),
    .B(_0590_),
    .X(_0606_));
 sky130_fd_sc_hd__inv_2 _1403_ (.A(_0594_),
    .Y(_0607_));
 sky130_fd_sc_hd__inv_2 _1404_ (.A(_0593_),
    .Y(_0608_));
 sky130_fd_sc_hd__o2bb2a_1 _1405_ (.A1_N(_0585_),
    .A2_N(_0586_),
    .B1(_0607_),
    .B2(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__and3_1 _1406_ (.A(_0605_),
    .B(_0606_),
    .C(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__a22o_1 _1407_ (.A1(_0607_),
    .A2(_0608_),
    .B1(_0592_),
    .B2(_0590_),
    .X(_0611_));
 sky130_fd_sc_hd__a21oi_1 _1408_ (.A1(_0603_),
    .A2(_0598_),
    .B1(_0604_),
    .Y(_0612_));
 sky130_fd_sc_hd__a31o_1 _1409_ (.A1(_0605_),
    .A2(_0611_),
    .A3(_0606_),
    .B1(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__a31o_1 _1410_ (.A1(_0588_),
    .A2(_0595_),
    .A3(_0610_),
    .B1(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _1411_ (.A0(\MAC.add.b1[8] ),
    .A1(\MAC.add.a1[8] ),
    .S(_0538_),
    .X(_0615_));
 sky130_fd_sc_hd__and4bb_1 _1412_ (.A_N(_0615_),
    .B_N(_0513_),
    .C(_0506_),
    .D(_0534_),
    .X(_0616_));
 sky130_fd_sc_hd__a31o_4 _1413_ (.A1(_0506_),
    .A2(_0567_),
    .A3(_0614_),
    .B1(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_2 _1414_ (.A0(_0565_),
    .A1(_0566_),
    .S(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _1415_ (.A0(\MAC.add.a1[0] ),
    .A1(\MAC.add.b1[0] ),
    .S(_0553_),
    .X(_0619_));
 sky130_fd_sc_hd__a31oi_1 _1416_ (.A1(_0506_),
    .A2(_0567_),
    .A3(_0614_),
    .B1(_0616_),
    .Y(_0620_));
 sky130_fd_sc_hd__a311o_1 _1417_ (.A1(_0506_),
    .A2(_0567_),
    .A3(_0614_),
    .B1(_0616_),
    .C1(_0549_),
    .X(_0621_));
 sky130_fd_sc_hd__xor2_4 _1418_ (.A(\MAC.add.a1[15] ),
    .B(\MAC.add.b1[15] ),
    .X(_0622_));
 sky130_fd_sc_hd__o211a_1 _1419_ (.A1(_0619_),
    .A2(_0620_),
    .B1(_0621_),
    .C1(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__xnor2_2 _1420_ (.A(_0618_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__clkbuf_4 _1421_ (.A(_0620_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _1422_ (.A0(_0565_),
    .A1(_0566_),
    .S(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__xnor2_2 _1423_ (.A(_0624_),
    .B(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__xnor2_2 _1424_ (.A(_0555_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__o21a_1 _1425_ (.A1(_0619_),
    .A2(_0625_),
    .B1(_0621_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_2 _1426_ (.A0(_0573_),
    .A1(_0574_),
    .S(_0617_),
    .X(_0630_));
 sky130_fd_sc_hd__inv_2 _1427_ (.A(_0585_),
    .Y(_0631_));
 sky130_fd_sc_hd__mux2_1 _1428_ (.A0(_0631_),
    .A1(_0586_),
    .S(_0617_),
    .X(_0632_));
 sky130_fd_sc_hd__or4_4 _1429_ (.A(_0629_),
    .B(_0618_),
    .C(_0630_),
    .D(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_2 _1430_ (.A0(_0607_),
    .A1(_0593_),
    .S(_0617_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _1431_ (.A0(_0592_),
    .A1(_0589_),
    .S(_0617_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _1432_ (.A0(_0600_),
    .A1(_0601_),
    .S(_0617_),
    .X(_0636_));
 sky130_fd_sc_hd__or4_4 _1433_ (.A(_0633_),
    .B(_0634_),
    .C(_0635_),
    .D(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_2 _1434_ (.A0(_0597_),
    .A1(_0598_),
    .S(_0617_),
    .X(_0638_));
 sky130_fd_sc_hd__nor2_1 _1435_ (.A(_0514_),
    .B(_0596_),
    .Y(_0639_));
 sky130_fd_sc_hd__o41a_1 _1436_ (.A1(_0506_),
    .A2(_0637_),
    .A3(_0638_),
    .A4(_0639_),
    .B1(_0622_),
    .X(_0640_));
 sky130_fd_sc_hd__o21ai_2 _1437_ (.A1(_0637_),
    .A2(_0638_),
    .B1(_0622_),
    .Y(_0641_));
 sky130_fd_sc_hd__mux2_1 _1438_ (.A0(_0615_),
    .A1(_0639_),
    .S(_0625_),
    .X(_0642_));
 sky130_fd_sc_hd__xnor2_2 _1439_ (.A(_0641_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__mux2_2 _1440_ (.A0(_0615_),
    .A1(_0639_),
    .S(_0617_),
    .X(_0644_));
 sky130_fd_sc_hd__nand2_1 _1441_ (.A(_0643_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__o31a_1 _1442_ (.A1(_0633_),
    .A2(_0634_),
    .A3(_0635_),
    .B1(_0622_),
    .X(_0646_));
 sky130_fd_sc_hd__xnor2_1 _1443_ (.A(_0636_),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(_0600_),
    .A1(_0601_),
    .S(_0625_),
    .X(_0648_));
 sky130_fd_sc_hd__inv_2 _1445_ (.A(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__nor2_2 _1446_ (.A(_0647_),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__and2_1 _1447_ (.A(_0647_),
    .B(_0649_),
    .X(_0651_));
 sky130_fd_sc_hd__nor2_1 _1448_ (.A(_0650_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__o21ai_1 _1449_ (.A1(_0633_),
    .A2(_0634_),
    .B1(_0622_),
    .Y(_0653_));
 sky130_fd_sc_hd__xnor2_1 _1450_ (.A(_0635_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(_0592_),
    .A1(_0589_),
    .S(_0625_),
    .X(_0655_));
 sky130_fd_sc_hd__or2_1 _1452_ (.A(_0654_),
    .B(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__xnor2_1 _1453_ (.A(\MAC.add.a1[15] ),
    .B(\MAC.add.b1[15] ),
    .Y(_0657_));
 sky130_fd_sc_hd__nor4_1 _1454_ (.A(_0629_),
    .B(_0618_),
    .C(_0630_),
    .D(_0632_),
    .Y(_0658_));
 sky130_fd_sc_hd__nor2_1 _1455_ (.A(_0657_),
    .B(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__xnor2_2 _1456_ (.A(_0634_),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__mux2_2 _1457_ (.A0(_0594_),
    .A1(_0608_),
    .S(_0625_),
    .X(_0661_));
 sky130_fd_sc_hd__nand2_1 _1458_ (.A(_0660_),
    .B(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__o31a_1 _1459_ (.A1(_0629_),
    .A2(_0618_),
    .A3(_0630_),
    .B1(_0622_),
    .X(_0663_));
 sky130_fd_sc_hd__xor2_1 _1460_ (.A(_0632_),
    .B(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _1461_ (.A0(_0631_),
    .A1(_0586_),
    .S(_0625_),
    .X(_0665_));
 sky130_fd_sc_hd__or2_2 _1462_ (.A(_0664_),
    .B(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__and2b_1 _1463_ (.A_N(_0624_),
    .B(_0626_),
    .X(_0667_));
 sky130_fd_sc_hd__a21o_1 _1464_ (.A1(_0555_),
    .A2(_0627_),
    .B1(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__o21a_1 _1465_ (.A1(_0629_),
    .A2(_0618_),
    .B1(_0622_),
    .X(_0669_));
 sky130_fd_sc_hd__xnor2_2 _1466_ (.A(_0630_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__inv_2 _1467_ (.A(_0573_),
    .Y(_0671_));
 sky130_fd_sc_hd__mux2_1 _1468_ (.A0(_0671_),
    .A1(_0575_),
    .S(_0625_),
    .X(_0672_));
 sky130_fd_sc_hd__inv_2 _1469_ (.A(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__xnor2_2 _1470_ (.A(_0670_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__and2_1 _1471_ (.A(_0664_),
    .B(_0665_),
    .X(_0675_));
 sky130_fd_sc_hd__nor2_1 _1472_ (.A(_0670_),
    .B(_0672_),
    .Y(_0676_));
 sky130_fd_sc_hd__a211o_1 _1473_ (.A1(_0668_),
    .A2(_0674_),
    .B1(_0675_),
    .C1(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__nor2_1 _1474_ (.A(_0660_),
    .B(_0661_),
    .Y(_0678_));
 sky130_fd_sc_hd__and2_1 _1475_ (.A(_0654_),
    .B(_0655_),
    .X(_0679_));
 sky130_fd_sc_hd__a311o_1 _1476_ (.A1(_0662_),
    .A2(_0666_),
    .A3(_0677_),
    .B1(_0678_),
    .C1(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(_0597_),
    .A1(_0598_),
    .S(_0625_),
    .X(_0681_));
 sky130_fd_sc_hd__nand2_1 _1478_ (.A(_0622_),
    .B(_0637_),
    .Y(_0682_));
 sky130_fd_sc_hd__xnor2_1 _1479_ (.A(_0638_),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__a32o_1 _1480_ (.A1(_0652_),
    .A2(_0656_),
    .A3(_0680_),
    .B1(_0681_),
    .B2(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__xor2_2 _1481_ (.A(_0643_),
    .B(_0644_),
    .X(_0685_));
 sky130_fd_sc_hd__or2_4 _1482_ (.A(_0683_),
    .B(_0681_),
    .X(_0686_));
 sky130_fd_sc_hd__o211ai_4 _1483_ (.A1(_0650_),
    .A2(_0684_),
    .B1(_0685_),
    .C1(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__o31a_1 _1484_ (.A1(_0637_),
    .A2(_0638_),
    .A3(_0642_),
    .B1(_0622_),
    .X(_0688_));
 sky130_fd_sc_hd__xnor2_2 _1485_ (.A(_0506_),
    .B(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__a31o_1 _1486_ (.A1(_0645_),
    .A2(_0687_),
    .A3(_0689_),
    .B1(_0457_),
    .X(_0690_));
 sky130_fd_sc_hd__or2_1 _1487_ (.A(_0640_),
    .B(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__buf_2 _1488_ (.A(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__a21oi_1 _1489_ (.A1(_0456_),
    .A2(_0625_),
    .B1(_0550_),
    .Y(_0693_));
 sky130_fd_sc_hd__a21oi_1 _1490_ (.A1(_0456_),
    .A2(_0617_),
    .B1(_0554_),
    .Y(_0694_));
 sky130_fd_sc_hd__nor2_1 _1491_ (.A(_0693_),
    .B(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__a31o_1 _1492_ (.A1(_0491_),
    .A2(_0549_),
    .A3(_0619_),
    .B1(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__a31o_1 _1493_ (.A1(_0652_),
    .A2(_0656_),
    .A3(_0680_),
    .B1(_0650_),
    .X(_0697_));
 sky130_fd_sc_hd__nand2_1 _1494_ (.A(_0683_),
    .B(_0681_),
    .Y(_0698_));
 sky130_fd_sc_hd__inv_2 _1495_ (.A(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__a211o_1 _1496_ (.A1(_0686_),
    .A2(_0697_),
    .B1(_0685_),
    .C1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__and2_1 _1497_ (.A(_0457_),
    .B(_0644_),
    .X(_0701_));
 sky130_fd_sc_hd__a31o_2 _1498_ (.A1(_0491_),
    .A2(_0687_),
    .A3(_0700_),
    .B1(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__a21oi_2 _1499_ (.A1(_0698_),
    .A2(_0686_),
    .B1(_0697_),
    .Y(_0703_));
 sky130_fd_sc_hd__a31o_1 _1500_ (.A1(_0698_),
    .A2(_0686_),
    .A3(_0697_),
    .B1(_0457_),
    .X(_0704_));
 sky130_fd_sc_hd__a31o_1 _1501_ (.A1(_0662_),
    .A2(_0666_),
    .A3(_0677_),
    .B1(_0678_),
    .X(_0705_));
 sky130_fd_sc_hd__or2b_1 _1502_ (.A(_0679_),
    .B_N(_0656_),
    .X(_0706_));
 sky130_fd_sc_hd__xor2_2 _1503_ (.A(_0705_),
    .B(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__xor2_1 _1504_ (.A(_0660_),
    .B(_0661_),
    .X(_0708_));
 sky130_fd_sc_hd__nand3_1 _1505_ (.A(_0708_),
    .B(_0666_),
    .C(_0677_),
    .Y(_0709_));
 sky130_fd_sc_hd__a21o_1 _1506_ (.A1(_0666_),
    .A2(_0677_),
    .B1(_0708_),
    .X(_0710_));
 sky130_fd_sc_hd__nor2_1 _1507_ (.A(_0491_),
    .B(_0661_),
    .Y(_0711_));
 sky130_fd_sc_hd__a31o_2 _1508_ (.A1(_0491_),
    .A2(_0709_),
    .A3(_0710_),
    .B1(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__xor2_1 _1509_ (.A(_0668_),
    .B(_0674_),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_2 _1510_ (.A0(_0673_),
    .A1(_0713_),
    .S(_0491_),
    .X(_0714_));
 sky130_fd_sc_hd__nand2_1 _1511_ (.A(_0456_),
    .B(_0626_),
    .Y(_0715_));
 sky130_fd_sc_hd__o21ai_2 _1512_ (.A1(_0456_),
    .A2(_0628_),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__nor2_1 _1513_ (.A(_0716_),
    .B(_0696_),
    .Y(_0717_));
 sky130_fd_sc_hd__nand2_1 _1514_ (.A(_0456_),
    .B(_0665_),
    .Y(_0718_));
 sky130_fd_sc_hd__inv_2 _1515_ (.A(_0666_),
    .Y(_0719_));
 sky130_fd_sc_hd__a21oi_1 _1516_ (.A1(_0668_),
    .A2(_0674_),
    .B1(_0676_),
    .Y(_0720_));
 sky130_fd_sc_hd__nand2_1 _1517_ (.A(_0664_),
    .B(_0665_),
    .Y(_0721_));
 sky130_fd_sc_hd__a221o_1 _1518_ (.A1(_0721_),
    .A2(_0666_),
    .B1(_0668_),
    .B2(_0674_),
    .C1(_0676_),
    .X(_0722_));
 sky130_fd_sc_hd__o311ai_2 _1519_ (.A1(_0675_),
    .A2(_0719_),
    .A3(_0720_),
    .B1(_0722_),
    .C1(_0491_),
    .Y(_0723_));
 sky130_fd_sc_hd__o211a_1 _1520_ (.A1(_0714_),
    .A2(_0717_),
    .B1(_0718_),
    .C1(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__nand2_1 _1521_ (.A(_0457_),
    .B(_0655_),
    .Y(_0725_));
 sky130_fd_sc_hd__o221a_1 _1522_ (.A1(_0457_),
    .A2(_0707_),
    .B1(_0712_),
    .B2(_0724_),
    .C1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__nand3_1 _1523_ (.A(_0652_),
    .B(_0656_),
    .C(_0680_),
    .Y(_0727_));
 sky130_fd_sc_hd__a21o_1 _1524_ (.A1(_0656_),
    .A2(_0680_),
    .B1(_0652_),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_1 _1525_ (.A(_0491_),
    .B(_0649_),
    .Y(_0729_));
 sky130_fd_sc_hd__a31o_2 _1526_ (.A1(_0491_),
    .A2(_0727_),
    .A3(_0728_),
    .B1(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__nand2_1 _1527_ (.A(_0457_),
    .B(_0681_),
    .Y(_0731_));
 sky130_fd_sc_hd__o221a_1 _1528_ (.A1(_0703_),
    .A2(_0704_),
    .B1(_0726_),
    .B2(_0730_),
    .C1(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__a31oi_2 _1529_ (.A1(_0645_),
    .A2(_0687_),
    .A3(_0689_),
    .B1(_0457_),
    .Y(_0733_));
 sky130_fd_sc_hd__a21o_1 _1530_ (.A1(_0645_),
    .A2(_0687_),
    .B1(_0689_),
    .X(_0734_));
 sky130_fd_sc_hd__o211a_4 _1531_ (.A1(_0702_),
    .A2(_0732_),
    .B1(_0733_),
    .C1(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__nor2_1 _1532_ (.A(_0696_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__nand2_1 _1533_ (.A(_0733_),
    .B(_0734_),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _1534_ (.A(_0718_),
    .B(_0723_),
    .Y(_0738_));
 sky130_fd_sc_hd__or2_1 _1535_ (.A(_0738_),
    .B(_0714_),
    .X(_0739_));
 sky130_fd_sc_hd__o21ai_2 _1536_ (.A1(_0457_),
    .A2(_0707_),
    .B1(_0725_),
    .Y(_0740_));
 sky130_fd_sc_hd__nor2_1 _1537_ (.A(_0740_),
    .B(_0712_),
    .Y(_0741_));
 sky130_fd_sc_hd__o21ai_4 _1538_ (.A1(_0703_),
    .A2(_0704_),
    .B1(_0731_),
    .Y(_0742_));
 sky130_fd_sc_hd__a211o_1 _1539_ (.A1(_0739_),
    .A2(_0741_),
    .B1(_0730_),
    .C1(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__or3b_1 _1540_ (.A(_0737_),
    .B(_0702_),
    .C_N(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__clkbuf_4 _1541_ (.A(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__or2_1 _1542_ (.A(_0739_),
    .B(_0712_),
    .X(_0746_));
 sky130_fd_sc_hd__nor2_1 _1543_ (.A(_0740_),
    .B(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__or3_1 _1544_ (.A(_0730_),
    .B(_0702_),
    .C(_0742_),
    .X(_0748_));
 sky130_fd_sc_hd__or3_2 _1545_ (.A(_0737_),
    .B(_0747_),
    .C(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__and3_1 _1546_ (.A(_0736_),
    .B(_0745_),
    .C(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__or3_1 _1547_ (.A(_0740_),
    .B(_0746_),
    .C(_0748_),
    .X(_0751_));
 sky130_fd_sc_hd__o21a_1 _1548_ (.A1(_0457_),
    .A2(_0628_),
    .B1(_0715_),
    .X(_0752_));
 sky130_fd_sc_hd__nand2_1 _1549_ (.A(_0752_),
    .B(_0696_),
    .Y(_0753_));
 sky130_fd_sc_hd__inv_2 _1550_ (.A(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__o31a_1 _1551_ (.A1(_0737_),
    .A2(_0751_),
    .A3(_0754_),
    .B1(_0692_),
    .X(_0755_));
 sky130_fd_sc_hd__nand2_1 _1552_ (.A(_0750_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__o31a_1 _1553_ (.A1(_0457_),
    .A2(_0628_),
    .A3(_0692_),
    .B1(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_2 _1554_ (.A0(\MAC.add.b1[13] ),
    .A1(\MAC.add.a1[13] ),
    .S(_0538_),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_1 _1555_ (.A0(\MAC.add.b1[12] ),
    .A1(\MAC.add.a1[12] ),
    .S(_0538_),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_2 _1556_ (.A0(\MAC.add.b1[9] ),
    .A1(\MAC.add.a1[9] ),
    .S(_0538_),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_2 _1557_ (.A0(\MAC.add.b1[10] ),
    .A1(\MAC.add.a1[10] ),
    .S(_0538_),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _1558_ (.A0(\MAC.add.b1[11] ),
    .A1(\MAC.add.a1[11] ),
    .S(_0538_),
    .X(_0762_));
 sky130_fd_sc_hd__nor3_1 _1559_ (.A(_0760_),
    .B(_0761_),
    .C(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__xor2_1 _1560_ (.A(_0759_),
    .B(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__or2_1 _1561_ (.A(_0702_),
    .B(_0742_),
    .X(_0765_));
 sky130_fd_sc_hd__or2_1 _1562_ (.A(_0716_),
    .B(_0696_),
    .X(_0766_));
 sky130_fd_sc_hd__nor2_1 _1563_ (.A(_0746_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__and3_1 _1564_ (.A(_0640_),
    .B(_0733_),
    .C(_0734_),
    .X(_0768_));
 sky130_fd_sc_hd__clkbuf_2 _1565_ (.A(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__o41a_1 _1566_ (.A1(_0740_),
    .A2(_0730_),
    .A3(_0765_),
    .A4(_0767_),
    .B1(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__or2_1 _1567_ (.A(_0770_),
    .B(_0762_),
    .X(_0771_));
 sky130_fd_sc_hd__nor2_2 _1568_ (.A(_0640_),
    .B(_0690_),
    .Y(_0772_));
 sky130_fd_sc_hd__or2_1 _1569_ (.A(_0772_),
    .B(_0735_),
    .X(_0773_));
 sky130_fd_sc_hd__nor2_1 _1570_ (.A(_0740_),
    .B(_0730_),
    .Y(_0774_));
 sky130_fd_sc_hd__nor2_1 _1571_ (.A(_0714_),
    .B(_0766_),
    .Y(_0775_));
 sky130_fd_sc_hd__or3_1 _1572_ (.A(_0738_),
    .B(_0712_),
    .C(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__a211o_1 _1573_ (.A1(_0774_),
    .A2(_0776_),
    .B1(_0702_),
    .C1(_0742_),
    .X(_0777_));
 sky130_fd_sc_hd__a21o_1 _1574_ (.A1(_0769_),
    .A2(_0777_),
    .B1(_0761_),
    .X(_0778_));
 sky130_fd_sc_hd__and3_1 _1575_ (.A(_0769_),
    .B(_0777_),
    .C(_0761_),
    .X(_0779_));
 sky130_fd_sc_hd__a31o_1 _1576_ (.A1(_0773_),
    .A2(_0760_),
    .A3(_0778_),
    .B1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__and2_1 _1577_ (.A(_0770_),
    .B(_0762_),
    .X(_0781_));
 sky130_fd_sc_hd__a21o_1 _1578_ (.A1(_0771_),
    .A2(_0780_),
    .B1(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__o21a_1 _1579_ (.A1(_0751_),
    .A2(_0716_),
    .B1(_0769_),
    .X(_0783_));
 sky130_fd_sc_hd__and2_1 _1580_ (.A(_0759_),
    .B(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__nor2_1 _1581_ (.A(\MAC.add.a1[14] ),
    .B(\MAC.add.b1[14] ),
    .Y(_0785_));
 sky130_fd_sc_hd__or3b_1 _1582_ (.A(_0758_),
    .B(_0759_),
    .C_N(_0763_),
    .X(_0786_));
 sky130_fd_sc_hd__xnor2_1 _1583_ (.A(_0785_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__or2_1 _1584_ (.A(_0783_),
    .B(_0764_),
    .X(_0788_));
 sky130_fd_sc_hd__o311a_1 _1585_ (.A1(_0782_),
    .A2(_0763_),
    .A3(_0784_),
    .B1(_0787_),
    .C1(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__o21a_1 _1586_ (.A1(_0751_),
    .A2(_0753_),
    .B1(_0769_),
    .X(_0790_));
 sky130_fd_sc_hd__nand2_1 _1587_ (.A(_0785_),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__or4_4 _1588_ (.A(_0758_),
    .B(_0764_),
    .C(_0789_),
    .D(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__and4_1 _1589_ (.A(\MAC.add.a1[10] ),
    .B(\MAC.add.a1[9] ),
    .C(\MAC.add.a1[15] ),
    .D(\MAC.add.a1[0] ),
    .X(_0793_));
 sky130_fd_sc_hd__and3_1 _1590_ (.A(\MAC.add.a1[14] ),
    .B(\MAC.add.a1[13] ),
    .C(\MAC.add.a1[12] ),
    .X(_0794_));
 sky130_fd_sc_hd__and3_1 _1591_ (.A(\MAC.add.a1[11] ),
    .B(_0793_),
    .C(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__and4_1 _1592_ (.A(\MAC.add.a1[1] ),
    .B(\MAC.add.a1[2] ),
    .C(\MAC.add.a1[3] ),
    .D(\MAC.add.a1[4] ),
    .X(_0796_));
 sky130_fd_sc_hd__and4_1 _1593_ (.A(\MAC.add.a1[5] ),
    .B(\MAC.add.a1[6] ),
    .C(\MAC.add.a1[7] ),
    .D(\MAC.add.a1[8] ),
    .X(_0797_));
 sky130_fd_sc_hd__and4_1 _1594_ (.A(\MAC.add.b1[10] ),
    .B(\MAC.add.b1[9] ),
    .C(\MAC.add.b1[15] ),
    .D(\MAC.add.b1[0] ),
    .X(_0798_));
 sky130_fd_sc_hd__and4_1 _1595_ (.A(\MAC.add.b1[14] ),
    .B(\MAC.add.b1[13] ),
    .C(\MAC.add.b1[12] ),
    .D(\MAC.add.b1[11] ),
    .X(_0799_));
 sky130_fd_sc_hd__and4_1 _1596_ (.A(\MAC.add.b1[5] ),
    .B(\MAC.add.b1[6] ),
    .C(\MAC.add.b1[7] ),
    .D(\MAC.add.b1[8] ),
    .X(_0800_));
 sky130_fd_sc_hd__and4_1 _1597_ (.A(\MAC.add.b1[1] ),
    .B(\MAC.add.b1[2] ),
    .C(\MAC.add.b1[3] ),
    .D(\MAC.add.b1[4] ),
    .X(_0801_));
 sky130_fd_sc_hd__and4_1 _1598_ (.A(_0798_),
    .B(_0799_),
    .C(_0800_),
    .D(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__a31oi_2 _1599_ (.A1(_0795_),
    .A2(_0796_),
    .A3(_0797_),
    .B1(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__nand2_1 _1600_ (.A(_0773_),
    .B(_0760_),
    .Y(_0804_));
 sky130_fd_sc_hd__nand2_1 _1601_ (.A(_0769_),
    .B(_0777_),
    .Y(_0805_));
 sky130_fd_sc_hd__and3_1 _1602_ (.A(_0761_),
    .B(_0759_),
    .C(_0762_),
    .X(_0806_));
 sky130_fd_sc_hd__and4bb_1 _1603_ (.A_N(_0785_),
    .B_N(_0770_),
    .C(_0758_),
    .D(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__and4bb_1 _1604_ (.A_N(_0790_),
    .B_N(_0804_),
    .C(_0805_),
    .D(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__clkbuf_2 _1605_ (.A(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__a31oi_1 _1606_ (.A1(_0757_),
    .A2(_0792_),
    .A3(_0803_),
    .B1(_0809_),
    .Y(\MAC.add.c_add[0] ));
 sky130_fd_sc_hd__a211o_1 _1607_ (.A1(_0747_),
    .A2(_0754_),
    .B1(_0748_),
    .C1(_0737_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _1608_ (.A0(_0752_),
    .A1(_0696_),
    .S(_0735_),
    .X(_0811_));
 sky130_fd_sc_hd__inv_2 _1609_ (.A(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__a31o_1 _1610_ (.A1(_0745_),
    .A2(_0810_),
    .A3(_0812_),
    .B1(_0772_),
    .X(_0813_));
 sky130_fd_sc_hd__or2_1 _1611_ (.A(_0714_),
    .B(_0692_),
    .X(_0814_));
 sky130_fd_sc_hd__or2b_1 _1612_ (.A(_0809_),
    .B_N(_0803_),
    .X(_0815_));
 sky130_fd_sc_hd__clkbuf_2 _1613_ (.A(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__a21o_1 _1614_ (.A1(_0813_),
    .A2(_0814_),
    .B1(_0816_),
    .X(\MAC.add.c_add[1] ));
 sky130_fd_sc_hd__mux2_1 _1615_ (.A0(_0714_),
    .A1(_0716_),
    .S(_0735_),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_1 _1616_ (.A0(_0736_),
    .A1(_0817_),
    .S(_0745_),
    .X(_0818_));
 sky130_fd_sc_hd__a21o_1 _1617_ (.A1(_0810_),
    .A2(_0818_),
    .B1(_0772_),
    .X(_0819_));
 sky130_fd_sc_hd__o21a_1 _1618_ (.A1(_0738_),
    .A2(_0692_),
    .B1(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__buf_4 _1619_ (.A(_0792_),
    .X(_0821_));
 sky130_fd_sc_hd__o21a_1 _1620_ (.A1(_0816_),
    .A2(_0820_),
    .B1(_0821_),
    .X(\MAC.add.c_add[2] ));
 sky130_fd_sc_hd__mux2_1 _1621_ (.A0(_0738_),
    .A1(_0714_),
    .S(_0735_),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _1622_ (.A0(_0812_),
    .A1(_0822_),
    .S(_0745_),
    .X(_0823_));
 sky130_fd_sc_hd__a21oi_1 _1623_ (.A1(_0810_),
    .A2(_0823_),
    .B1(_0772_),
    .Y(_0824_));
 sky130_fd_sc_hd__o21ba_1 _1624_ (.A1(_0712_),
    .A2(_0692_),
    .B1_N(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__o21a_1 _1625_ (.A1(_0816_),
    .A2(_0825_),
    .B1(_0821_),
    .X(\MAC.add.c_add[3] ));
 sky130_fd_sc_hd__inv_2 _1626_ (.A(_0749_),
    .Y(_0826_));
 sky130_fd_sc_hd__mux2_1 _1627_ (.A0(_0712_),
    .A1(_0738_),
    .S(_0735_),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_1 _1628_ (.A0(_0817_),
    .A1(_0827_),
    .S(_0745_),
    .X(_0828_));
 sky130_fd_sc_hd__or2_1 _1629_ (.A(_0826_),
    .B(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__a21o_1 _1630_ (.A1(_0736_),
    .A2(_0745_),
    .B1(_0749_),
    .X(_0830_));
 sky130_fd_sc_hd__a31oi_2 _1631_ (.A1(_0795_),
    .A2(_0796_),
    .A3(_0797_),
    .B1(_0802_),
    .Y(_0831_));
 sky130_fd_sc_hd__o21ai_1 _1632_ (.A1(_0707_),
    .A2(_0692_),
    .B1(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__a311o_1 _1633_ (.A1(_0692_),
    .A2(_0829_),
    .A3(_0830_),
    .B1(_0832_),
    .C1(_0809_),
    .X(_0833_));
 sky130_fd_sc_hd__and2_1 _1634_ (.A(_0792_),
    .B(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__clkbuf_1 _1635_ (.A(_0834_),
    .X(\MAC.add.c_add[4] ));
 sky130_fd_sc_hd__or4_1 _1636_ (.A(\MAC.add.a1[14] ),
    .B(\MAC.add.b1[14] ),
    .C(_0758_),
    .D(_0764_),
    .X(_0835_));
 sky130_fd_sc_hd__or3b_1 _1637_ (.A(_0789_),
    .B(_0835_),
    .C_N(_0790_),
    .X(_0836_));
 sky130_fd_sc_hd__inv_2 _1638_ (.A(_0831_),
    .Y(_0837_));
 sky130_fd_sc_hd__inv_2 _1639_ (.A(_0745_),
    .Y(_0838_));
 sky130_fd_sc_hd__nor2_1 _1640_ (.A(_0838_),
    .B(_0811_),
    .Y(_0839_));
 sky130_fd_sc_hd__mux2_1 _1641_ (.A0(_0740_),
    .A1(_0712_),
    .S(_0735_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _1642_ (.A0(_0822_),
    .A1(_0840_),
    .S(_0745_),
    .X(_0841_));
 sky130_fd_sc_hd__o211a_1 _1643_ (.A1(_0749_),
    .A2(_0839_),
    .B1(_0841_),
    .C1(_0755_),
    .X(_0842_));
 sky130_fd_sc_hd__a211o_1 _1644_ (.A1(_0730_),
    .A2(_0772_),
    .B1(_0837_),
    .C1(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__a21o_1 _1645_ (.A1(_0836_),
    .A2(_0843_),
    .B1(_0809_),
    .X(\MAC.add.c_add[5] ));
 sky130_fd_sc_hd__mux2_1 _1646_ (.A0(_0730_),
    .A1(_0740_),
    .S(_0735_),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_1 _1647_ (.A0(_0827_),
    .A1(_0844_),
    .S(_0745_),
    .X(_0845_));
 sky130_fd_sc_hd__or2_1 _1648_ (.A(_0749_),
    .B(_0818_),
    .X(_0846_));
 sky130_fd_sc_hd__o211a_1 _1649_ (.A1(_0826_),
    .A2(_0845_),
    .B1(_0846_),
    .C1(_0755_),
    .X(_0847_));
 sky130_fd_sc_hd__a211o_1 _1650_ (.A1(_0742_),
    .A2(_0772_),
    .B1(_0837_),
    .C1(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__a21o_1 _1651_ (.A1(_0836_),
    .A2(_0848_),
    .B1(_0809_),
    .X(\MAC.add.c_add[6] ));
 sky130_fd_sc_hd__mux2_1 _1652_ (.A0(_0742_),
    .A1(_0730_),
    .S(_0735_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _1653_ (.A0(_0840_),
    .A1(_0849_),
    .S(_0745_),
    .X(_0850_));
 sky130_fd_sc_hd__a211o_1 _1654_ (.A1(_0826_),
    .A2(_0823_),
    .B1(_0850_),
    .C1(_0772_),
    .X(_0851_));
 sky130_fd_sc_hd__o21a_1 _1655_ (.A1(_0702_),
    .A2(_0692_),
    .B1(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__o21a_1 _1656_ (.A1(_0816_),
    .A2(_0852_),
    .B1(_0821_),
    .X(\MAC.add.c_add[7] ));
 sky130_fd_sc_hd__nor2_1 _1657_ (.A(_0750_),
    .B(_0828_),
    .Y(_0853_));
 sky130_fd_sc_hd__o21ai_1 _1658_ (.A1(_0737_),
    .A2(_0742_),
    .B1(_0702_),
    .Y(_0854_));
 sky130_fd_sc_hd__nand2_1 _1659_ (.A(_0838_),
    .B(_0844_),
    .Y(_0855_));
 sky130_fd_sc_hd__o2111a_1 _1660_ (.A1(_0810_),
    .A2(_0853_),
    .B1(_0854_),
    .C1(_0855_),
    .D1(_0692_),
    .X(_0856_));
 sky130_fd_sc_hd__a21oi_1 _1661_ (.A1(_0734_),
    .A2(_0772_),
    .B1(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__o21a_1 _1662_ (.A1(_0816_),
    .A2(_0857_),
    .B1(_0821_),
    .X(\MAC.add.c_add[8] ));
 sky130_fd_sc_hd__or2_1 _1663_ (.A(_0773_),
    .B(_0760_),
    .X(_0858_));
 sky130_fd_sc_hd__nand2_1 _1664_ (.A(_0804_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__a31oi_1 _1665_ (.A1(_0821_),
    .A2(_0803_),
    .A3(_0859_),
    .B1(_0809_),
    .Y(\MAC.add.c_add[9] ));
 sky130_fd_sc_hd__a21oi_1 _1666_ (.A1(_0769_),
    .A2(_0777_),
    .B1(_0761_),
    .Y(_0860_));
 sky130_fd_sc_hd__nor2_1 _1667_ (.A(_0860_),
    .B(_0779_),
    .Y(_0861_));
 sky130_fd_sc_hd__xnor2_1 _1668_ (.A(_0804_),
    .B(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__o31a_1 _1669_ (.A1(_0809_),
    .A2(_0837_),
    .A3(_0862_),
    .B1(_0821_),
    .X(\MAC.add.c_add[10] ));
 sky130_fd_sc_hd__or2b_1 _1670_ (.A(_0781_),
    .B_N(_0771_),
    .X(_0863_));
 sky130_fd_sc_hd__xnor2_1 _1671_ (.A(_0863_),
    .B(_0780_),
    .Y(_0864_));
 sky130_fd_sc_hd__o21a_1 _1672_ (.A1(_0816_),
    .A2(_0864_),
    .B1(_0821_),
    .X(\MAC.add.c_add[11] ));
 sky130_fd_sc_hd__or2_1 _1673_ (.A(_0759_),
    .B(_0783_),
    .X(_0865_));
 sky130_fd_sc_hd__or2b_1 _1674_ (.A(_0784_),
    .B_N(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__xnor2_1 _1675_ (.A(_0782_),
    .B(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__o21a_1 _1676_ (.A1(_0816_),
    .A2(_0867_),
    .B1(_0821_),
    .X(\MAC.add.c_add[12] ));
 sky130_fd_sc_hd__xnor2_1 _1677_ (.A(_0790_),
    .B(_0758_),
    .Y(_0868_));
 sky130_fd_sc_hd__a21oi_1 _1678_ (.A1(_0782_),
    .A2(_0865_),
    .B1(_0784_),
    .Y(_0869_));
 sky130_fd_sc_hd__xor2_1 _1679_ (.A(_0868_),
    .B(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__o21a_1 _1680_ (.A1(_0816_),
    .A2(_0870_),
    .B1(_0821_),
    .X(\MAC.add.c_add[13] ));
 sky130_fd_sc_hd__nand2_1 _1681_ (.A(_0790_),
    .B(_0758_),
    .Y(_0871_));
 sky130_fd_sc_hd__o21a_1 _1682_ (.A1(_0868_),
    .A2(_0869_),
    .B1(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__or2_1 _1683_ (.A(_0785_),
    .B(_0790_),
    .X(_0873_));
 sky130_fd_sc_hd__and2_1 _1684_ (.A(_0791_),
    .B(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__inv_2 _1685_ (.A(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__nor2_1 _1686_ (.A(_0872_),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__and2_1 _1687_ (.A(_0872_),
    .B(_0875_),
    .X(_0877_));
 sky130_fd_sc_hd__o31a_1 _1688_ (.A1(_0816_),
    .A2(_0876_),
    .A3(_0877_),
    .B1(_0821_),
    .X(\MAC.add.c_add[14] ));
 sky130_fd_sc_hd__or2_1 _1689_ (.A(\MAC.a[14] ),
    .B(\MAC.b[14] ),
    .X(_0878_));
 sky130_fd_sc_hd__and2_1 _1690_ (.A(\MAC.a[12] ),
    .B(\MAC.b[12] ),
    .X(_0879_));
 sky130_fd_sc_hd__nor2_1 _1691_ (.A(\MAC.a[12] ),
    .B(\MAC.b[12] ),
    .Y(_0880_));
 sky130_fd_sc_hd__or2_1 _1692_ (.A(_0879_),
    .B(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__nand2_1 _1693_ (.A(\MAC.a[10] ),
    .B(\MAC.b[10] ),
    .Y(_0882_));
 sky130_fd_sc_hd__or2_1 _1694_ (.A(\MAC.a[10] ),
    .B(\MAC.b[10] ),
    .X(_0883_));
 sky130_fd_sc_hd__nand2_1 _1695_ (.A(_0882_),
    .B(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__nand2_1 _1696_ (.A(\MAC.a[9] ),
    .B(\MAC.b[9] ),
    .Y(_0885_));
 sky130_fd_sc_hd__or2_1 _1697_ (.A(_0884_),
    .B(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__xnor2_1 _1698_ (.A(\MAC.a[11] ),
    .B(\MAC.b[11] ),
    .Y(_0887_));
 sky130_fd_sc_hd__a21oi_1 _1699_ (.A1(_0882_),
    .A2(_0886_),
    .B1(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__a21oi_1 _1700_ (.A1(\MAC.a[11] ),
    .A2(\MAC.b[11] ),
    .B1(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_1 _1701_ (.A(_0881_),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__xor2_1 _1702_ (.A(\MAC.a[13] ),
    .B(\MAC.b[13] ),
    .X(_0891_));
 sky130_fd_sc_hd__o21a_1 _1703_ (.A1(_0879_),
    .A2(_0890_),
    .B1(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__a21o_1 _1704_ (.A1(\MAC.a[13] ),
    .A2(\MAC.b[13] ),
    .B1(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__nand2_1 _1705_ (.A(\MAC.a[14] ),
    .B(\MAC.b[14] ),
    .Y(_0894_));
 sky130_fd_sc_hd__a21bo_1 _1706_ (.A1(_0878_),
    .A2(_0893_),
    .B1_N(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__nand2_1 _1707_ (.A(_0894_),
    .B(_0878_),
    .Y(_0896_));
 sky130_fd_sc_hd__xor2_1 _1708_ (.A(_0896_),
    .B(_0893_),
    .X(_0897_));
 sky130_fd_sc_hd__nor3_1 _1709_ (.A(_0879_),
    .B(_0890_),
    .C(_0891_),
    .Y(_0898_));
 sky130_fd_sc_hd__or2_1 _1710_ (.A(_0892_),
    .B(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__and2_1 _1711_ (.A(_0881_),
    .B(_0889_),
    .X(_0900_));
 sky130_fd_sc_hd__or2_1 _1712_ (.A(_0890_),
    .B(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__or2_1 _1713_ (.A(\MAC.a[9] ),
    .B(\MAC.b[9] ),
    .X(_0902_));
 sky130_fd_sc_hd__nand2_1 _1714_ (.A(_0885_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__or2_1 _1715_ (.A(_0884_),
    .B(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__and3_1 _1716_ (.A(_0882_),
    .B(_0886_),
    .C(_0887_),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_1 _1717_ (.A(_0888_),
    .B(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__xor2_1 _1718_ (.A(_0904_),
    .B(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__nand2_1 _1719_ (.A(_0884_),
    .B(_0885_),
    .Y(_0908_));
 sky130_fd_sc_hd__and2_1 _1720_ (.A(_0886_),
    .B(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__nand2_1 _1721_ (.A(_0903_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__nor4_1 _1722_ (.A(_0899_),
    .B(_0901_),
    .C(_0907_),
    .D(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__buf_2 _1723_ (.A(\MAC.a[5] ),
    .X(_0912_));
 sky130_fd_sc_hd__buf_2 _1724_ (.A(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__buf_2 _1725_ (.A(\MAC.a[6] ),
    .X(_0914_));
 sky130_fd_sc_hd__buf_2 _1726_ (.A(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__and4_1 _1727_ (.A(\MAC.a[10] ),
    .B(\MAC.a[9] ),
    .C(\MAC.a[12] ),
    .D(\MAC.a[11] ),
    .X(_0916_));
 sky130_fd_sc_hd__and2_1 _1728_ (.A(\MAC.a[0] ),
    .B(\MAC.a[1] ),
    .X(_0917_));
 sky130_fd_sc_hd__and4_1 _1729_ (.A(_0913_),
    .B(_0915_),
    .C(_0916_),
    .D(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__buf_2 _1730_ (.A(\MAC.a[4] ),
    .X(_0919_));
 sky130_fd_sc_hd__buf_2 _1731_ (.A(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__buf_2 _1732_ (.A(\MAC.a[7] ),
    .X(_0921_));
 sky130_fd_sc_hd__buf_2 _1733_ (.A(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__buf_2 _1734_ (.A(\MAC.a[8] ),
    .X(_0923_));
 sky130_fd_sc_hd__buf_2 _1735_ (.A(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__and4_1 _1736_ (.A(_0920_),
    .B(_0922_),
    .C(_0924_),
    .D(\MAC.a[15] ),
    .X(_0925_));
 sky130_fd_sc_hd__buf_2 _1737_ (.A(\MAC.a[2] ),
    .X(_0926_));
 sky130_fd_sc_hd__buf_2 _1738_ (.A(\MAC.a[3] ),
    .X(_0927_));
 sky130_fd_sc_hd__buf_2 _1739_ (.A(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__and4_1 _1740_ (.A(\MAC.a[14] ),
    .B(\MAC.a[13] ),
    .C(_0926_),
    .D(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__buf_2 _1741_ (.A(\MAC.b[0] ),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_2 _1742_ (.A(\MAC.b[1] ),
    .X(_0931_));
 sky130_fd_sc_hd__buf_2 _1743_ (.A(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__and4_1 _1744_ (.A(\MAC.b[10] ),
    .B(\MAC.b[9] ),
    .C(_0930_),
    .D(_0932_),
    .X(_0933_));
 sky130_fd_sc_hd__clkbuf_2 _1745_ (.A(\MAC.b[3] ),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_4 _1746_ (.A(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__clkbuf_2 _1747_ (.A(\MAC.b[4] ),
    .X(_0936_));
 sky130_fd_sc_hd__clkbuf_4 _1748_ (.A(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__buf_2 _1749_ (.A(\MAC.b[7] ),
    .X(_0938_));
 sky130_fd_sc_hd__buf_2 _1750_ (.A(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__buf_2 _1751_ (.A(\MAC.b[8] ),
    .X(_0940_));
 sky130_fd_sc_hd__buf_2 _1752_ (.A(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__and4_1 _1753_ (.A(_0935_),
    .B(_0937_),
    .C(_0939_),
    .D(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__and4_1 _1754_ (.A(\MAC.b[12] ),
    .B(\MAC.b[11] ),
    .C(\MAC.b[14] ),
    .D(\MAC.b[13] ),
    .X(_0943_));
 sky130_fd_sc_hd__clkbuf_2 _1755_ (.A(\MAC.b[2] ),
    .X(_0944_));
 sky130_fd_sc_hd__clkbuf_4 _1756_ (.A(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__clkbuf_2 _1757_ (.A(\MAC.b[5] ),
    .X(_0946_));
 sky130_fd_sc_hd__buf_2 _1758_ (.A(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__buf_2 _1759_ (.A(\MAC.b[6] ),
    .X(_0948_));
 sky130_fd_sc_hd__and4_1 _1760_ (.A(_0945_),
    .B(_0947_),
    .C(_0948_),
    .D(\MAC.b[15] ),
    .X(_0949_));
 sky130_fd_sc_hd__and4_1 _1761_ (.A(_0933_),
    .B(_0942_),
    .C(_0943_),
    .D(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__a31o_1 _1762_ (.A1(_0918_),
    .A2(_0925_),
    .A3(_0929_),
    .B1(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__a31oi_2 _1763_ (.A1(_0895_),
    .A2(_0897_),
    .A3(_0911_),
    .B1(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__and3_1 _1764_ (.A(_0915_),
    .B(_0922_),
    .C(_0941_),
    .X(_0953_));
 sky130_fd_sc_hd__a21oi_1 _1765_ (.A1(_0922_),
    .A2(_0941_),
    .B1(_0915_),
    .Y(_0954_));
 sky130_fd_sc_hd__and4bb_1 _1766_ (.A_N(_0953_),
    .B_N(_0954_),
    .C(_0924_),
    .D(_0939_),
    .X(_0955_));
 sky130_fd_sc_hd__nor2_1 _1767_ (.A(_0953_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__and2_1 _1768_ (.A(_0924_),
    .B(_0941_),
    .X(_0957_));
 sky130_fd_sc_hd__or2_1 _1769_ (.A(_0922_),
    .B(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__nand2_1 _1770_ (.A(_0922_),
    .B(_0957_),
    .Y(_0959_));
 sky130_fd_sc_hd__and3_1 _1771_ (.A(_0939_),
    .B(_0958_),
    .C(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__a21oi_1 _1772_ (.A1(_0958_),
    .A2(_0959_),
    .B1(_0939_),
    .Y(_0961_));
 sky130_fd_sc_hd__or3_1 _1773_ (.A(_0956_),
    .B(_0960_),
    .C(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__nand2_1 _1774_ (.A(_0921_),
    .B(_0938_),
    .Y(_0963_));
 sky130_fd_sc_hd__nor2_1 _1775_ (.A(_0924_),
    .B(_0941_),
    .Y(_0964_));
 sky130_fd_sc_hd__or3_1 _1776_ (.A(_0963_),
    .B(_0957_),
    .C(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__o21ai_1 _1777_ (.A1(_0957_),
    .A2(_0964_),
    .B1(_0959_),
    .Y(_0966_));
 sky130_fd_sc_hd__or2_1 _1778_ (.A(_0960_),
    .B(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__o21ai_1 _1779_ (.A1(_0960_),
    .A2(_0961_),
    .B1(_0956_),
    .Y(_0968_));
 sky130_fd_sc_hd__nand3_1 _1780_ (.A(_0913_),
    .B(_0915_),
    .C(_0941_),
    .Y(_0969_));
 sky130_fd_sc_hd__and3_1 _1781_ (.A(_0912_),
    .B(_0914_),
    .C(_0940_),
    .X(_0970_));
 sky130_fd_sc_hd__a21oi_1 _1782_ (.A1(_0915_),
    .A2(_0940_),
    .B1(_0913_),
    .Y(_0971_));
 sky130_fd_sc_hd__or3_1 _1783_ (.A(_0970_),
    .B(_0963_),
    .C(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__o2bb2a_1 _1784_ (.A1_N(_0924_),
    .A2_N(_0939_),
    .B1(_0953_),
    .B2(_0954_),
    .X(_0973_));
 sky130_fd_sc_hd__a211oi_1 _1785_ (.A1(_0969_),
    .A2(_0972_),
    .B1(_0955_),
    .C1(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__o211a_1 _1786_ (.A1(_0955_),
    .A2(_0973_),
    .B1(_0969_),
    .C1(_0972_),
    .X(_0975_));
 sky130_fd_sc_hd__nor2_1 _1787_ (.A(_0974_),
    .B(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__and3_1 _1788_ (.A(_0923_),
    .B(_0937_),
    .C(_0947_),
    .X(_0977_));
 sky130_fd_sc_hd__clkbuf_2 _1789_ (.A(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__a21o_1 _1790_ (.A1(_0976_),
    .A2(_0978_),
    .B1(_0974_),
    .X(_0979_));
 sky130_fd_sc_hd__and3_1 _1791_ (.A(_0962_),
    .B(_0968_),
    .C(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__and4_1 _1792_ (.A(_0962_),
    .B(_0965_),
    .C(_0967_),
    .D(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__nand2_1 _1793_ (.A(_0924_),
    .B(_0937_),
    .Y(_0982_));
 sky130_fd_sc_hd__a21oi_1 _1794_ (.A1(_0923_),
    .A2(_0947_),
    .B1(_0937_),
    .Y(_0983_));
 sky130_fd_sc_hd__nor2_1 _1795_ (.A(_0978_),
    .B(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__a22o_1 _1796_ (.A1(_0923_),
    .A2(_0937_),
    .B1(_0947_),
    .B2(_0921_),
    .X(_0985_));
 sky130_fd_sc_hd__nand2_1 _1797_ (.A(_0921_),
    .B(_0978_),
    .Y(_0986_));
 sky130_fd_sc_hd__and4_1 _1798_ (.A(_0935_),
    .B(_0984_),
    .C(_0985_),
    .D(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__and3_1 _1799_ (.A(_0947_),
    .B(_0982_),
    .C(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__and3_1 _1800_ (.A(_0920_),
    .B(_0913_),
    .C(_0941_),
    .X(_0989_));
 sky130_fd_sc_hd__nand3_1 _1801_ (.A(_0920_),
    .B(_0913_),
    .C(_0941_),
    .Y(_0990_));
 sky130_fd_sc_hd__a21o_1 _1802_ (.A1(_0913_),
    .A2(_0940_),
    .B1(_0920_),
    .X(_0991_));
 sky130_fd_sc_hd__and4_1 _1803_ (.A(_0915_),
    .B(_0939_),
    .C(_0990_),
    .D(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__o21ai_1 _1804_ (.A1(_0970_),
    .A2(_0971_),
    .B1(_0963_),
    .Y(_0993_));
 sky130_fd_sc_hd__o211a_1 _1805_ (.A1(_0989_),
    .A2(_0992_),
    .B1(_0972_),
    .C1(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__inv_2 _1806_ (.A(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__a211o_1 _1807_ (.A1(_0972_),
    .A2(_0993_),
    .B1(_0989_),
    .C1(_0992_),
    .X(_0996_));
 sky130_fd_sc_hd__and2_1 _1808_ (.A(_0995_),
    .B(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__a21oi_1 _1809_ (.A1(_0947_),
    .A2(_0982_),
    .B1(_0987_),
    .Y(_0998_));
 sky130_fd_sc_hd__nor2_1 _1810_ (.A(_0988_),
    .B(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__and2_1 _1811_ (.A(_0997_),
    .B(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__xor2_1 _1812_ (.A(_0976_),
    .B(_0978_),
    .X(_1001_));
 sky130_fd_sc_hd__o21a_1 _1813_ (.A1(_0988_),
    .A2(_1000_),
    .B1(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__nor3_1 _1814_ (.A(_1001_),
    .B(_0988_),
    .C(_1000_),
    .Y(_1003_));
 sky130_fd_sc_hd__or2_1 _1815_ (.A(_1002_),
    .B(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__nor2_1 _1816_ (.A(_0995_),
    .B(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__nand2_1 _1817_ (.A(_0962_),
    .B(_0968_),
    .Y(_1006_));
 sky130_fd_sc_hd__xnor2_1 _1818_ (.A(_1006_),
    .B(_0979_),
    .Y(_1007_));
 sky130_fd_sc_hd__o21ai_1 _1819_ (.A1(_1002_),
    .A2(_1005_),
    .B1(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__a31o_1 _1820_ (.A1(_0962_),
    .A2(_0965_),
    .A3(_0967_),
    .B1(_0980_),
    .X(_1009_));
 sky130_fd_sc_hd__or2b_1 _1821_ (.A(_0981_),
    .B_N(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__or2_1 _1822_ (.A(_1008_),
    .B(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_1 _1823_ (.A(_1008_),
    .B(_1010_),
    .Y(_1012_));
 sky130_fd_sc_hd__nand2_1 _1824_ (.A(_1011_),
    .B(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__nor2_1 _1825_ (.A(_0997_),
    .B(_0999_),
    .Y(_1014_));
 sky130_fd_sc_hd__or2_1 _1826_ (.A(_1000_),
    .B(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__a22oi_1 _1827_ (.A1(_0915_),
    .A2(_0939_),
    .B1(_0990_),
    .B2(_0991_),
    .Y(_1016_));
 sky130_fd_sc_hd__nor2_1 _1828_ (.A(_0992_),
    .B(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__and3_1 _1829_ (.A(_0928_),
    .B(_0920_),
    .C(_0940_),
    .X(_1018_));
 sky130_fd_sc_hd__a21o_1 _1830_ (.A1(_0919_),
    .A2(_0940_),
    .B1(_0928_),
    .X(_1019_));
 sky130_fd_sc_hd__and4b_1 _1831_ (.A_N(_1018_),
    .B(_1019_),
    .C(_0912_),
    .D(_0938_),
    .X(_1020_));
 sky130_fd_sc_hd__or2_1 _1832_ (.A(_1018_),
    .B(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__xnor2_1 _1833_ (.A(_1017_),
    .B(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__nand4_2 _1834_ (.A(_0914_),
    .B(_0921_),
    .C(_0937_),
    .D(_0947_),
    .Y(_1023_));
 sky130_fd_sc_hd__a22o_1 _1835_ (.A1(_0921_),
    .A2(_0937_),
    .B1(_0947_),
    .B2(_0914_),
    .X(_1024_));
 sky130_fd_sc_hd__nand4_1 _1836_ (.A(_0923_),
    .B(_0935_),
    .C(_1023_),
    .D(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__nand2_1 _1837_ (.A(_0985_),
    .B(_0986_),
    .Y(_1026_));
 sky130_fd_sc_hd__xor2_1 _1838_ (.A(_0935_),
    .B(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__a21oi_1 _1839_ (.A1(_1023_),
    .A2(_1025_),
    .B1(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__a221oi_1 _1840_ (.A1(_0922_),
    .A2(_0978_),
    .B1(_0985_),
    .B2(_0935_),
    .C1(_0984_),
    .Y(_1029_));
 sky130_fd_sc_hd__or3_1 _1841_ (.A(_0987_),
    .B(_1028_),
    .C(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__o21bai_1 _1842_ (.A1(_1022_),
    .A2(_1030_),
    .B1_N(_1028_),
    .Y(_1031_));
 sky130_fd_sc_hd__or2b_1 _1843_ (.A(_1015_),
    .B_N(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__or2b_1 _1844_ (.A(_1031_),
    .B_N(_1015_),
    .X(_1033_));
 sky130_fd_sc_hd__nand2_1 _1845_ (.A(_1032_),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__or4b_1 _1846_ (.A(_0992_),
    .B(_1016_),
    .C(_1034_),
    .D_N(_1021_),
    .X(_1035_));
 sky130_fd_sc_hd__and2_1 _1847_ (.A(_0995_),
    .B(_1004_),
    .X(_1036_));
 sky130_fd_sc_hd__or2_1 _1848_ (.A(_1005_),
    .B(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__a21oi_1 _1849_ (.A1(_1032_),
    .A2(_1035_),
    .B1(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__and3_1 _1850_ (.A(_1037_),
    .B(_1032_),
    .C(_1035_),
    .X(_1039_));
 sky130_fd_sc_hd__nor2_1 _1851_ (.A(_1038_),
    .B(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__and2_1 _1852_ (.A(_0948_),
    .B(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__or3_1 _1853_ (.A(_1002_),
    .B(_1005_),
    .C(_1007_),
    .X(_1042_));
 sky130_fd_sc_hd__and2_1 _1854_ (.A(_1008_),
    .B(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__o21a_1 _1855_ (.A1(_1038_),
    .A2(_1041_),
    .B1(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__nor2_1 _1856_ (.A(_0948_),
    .B(_1040_),
    .Y(_1045_));
 sky130_fd_sc_hd__or2_1 _1857_ (.A(_1041_),
    .B(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__xnor2_1 _1858_ (.A(_1022_),
    .B(_1030_),
    .Y(_1047_));
 sky130_fd_sc_hd__inv_2 _1859_ (.A(_1019_),
    .Y(_1048_));
 sky130_fd_sc_hd__o2bb2a_1 _1860_ (.A1_N(_0913_),
    .A2_N(_0938_),
    .B1(_1018_),
    .B2(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__nor2_1 _1861_ (.A(_1020_),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__and3_1 _1862_ (.A(_0926_),
    .B(_0928_),
    .C(_0940_),
    .X(_1051_));
 sky130_fd_sc_hd__a21o_1 _1863_ (.A1(_0927_),
    .A2(_0940_),
    .B1(_0926_),
    .X(_1052_));
 sky130_fd_sc_hd__and4b_1 _1864_ (.A_N(_1051_),
    .B(_1052_),
    .C(_0920_),
    .D(_0938_),
    .X(_1053_));
 sky130_fd_sc_hd__or2_1 _1865_ (.A(_1051_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__xor2_1 _1866_ (.A(_1050_),
    .B(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__and3_1 _1867_ (.A(_1027_),
    .B(_1023_),
    .C(_1025_),
    .X(_1056_));
 sky130_fd_sc_hd__or2_1 _1868_ (.A(_1028_),
    .B(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__a22o_1 _1869_ (.A1(_0923_),
    .A2(_0934_),
    .B1(_1023_),
    .B2(_1024_),
    .X(_1058_));
 sky130_fd_sc_hd__and2_1 _1870_ (.A(_1025_),
    .B(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__and4_1 _1871_ (.A(\MAC.a[5] ),
    .B(\MAC.a[6] ),
    .C(_0936_),
    .D(_0946_),
    .X(_1060_));
 sky130_fd_sc_hd__a22oi_1 _1872_ (.A1(\MAC.a[6] ),
    .A2(_0936_),
    .B1(_0947_),
    .B2(_0912_),
    .Y(_1061_));
 sky130_fd_sc_hd__and4bb_1 _1873_ (.A_N(_1060_),
    .B_N(_1061_),
    .C(_0921_),
    .D(_0934_),
    .X(_1062_));
 sky130_fd_sc_hd__nor2_1 _1874_ (.A(_1060_),
    .B(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__xnor2_1 _1875_ (.A(_1059_),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__and2b_1 _1876_ (.A_N(_1063_),
    .B(_1059_),
    .X(_1065_));
 sky130_fd_sc_hd__a21oi_1 _1877_ (.A1(_0945_),
    .A2(_1064_),
    .B1(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__xnor2_1 _1878_ (.A(_1057_),
    .B(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__inv_2 _1879_ (.A(_1067_),
    .Y(_1068_));
 sky130_fd_sc_hd__nor2_1 _1880_ (.A(_1057_),
    .B(_1066_),
    .Y(_1069_));
 sky130_fd_sc_hd__a21oi_1 _1881_ (.A1(_1055_),
    .A2(_1068_),
    .B1(_1069_),
    .Y(_1070_));
 sky130_fd_sc_hd__nor2_1 _1882_ (.A(_1047_),
    .B(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__and2_1 _1883_ (.A(_1050_),
    .B(_1054_),
    .X(_1072_));
 sky130_fd_sc_hd__inv_2 _1884_ (.A(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__xnor2_1 _1885_ (.A(_1047_),
    .B(_1070_),
    .Y(_1074_));
 sky130_fd_sc_hd__nor2_1 _1886_ (.A(_1073_),
    .B(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__and2_1 _1887_ (.A(_1017_),
    .B(_1021_),
    .X(_1076_));
 sky130_fd_sc_hd__xnor2_1 _1888_ (.A(_1076_),
    .B(_1034_),
    .Y(_1077_));
 sky130_fd_sc_hd__o21a_1 _1889_ (.A1(_1071_),
    .A2(_1075_),
    .B1(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__nor3_1 _1890_ (.A(_1077_),
    .B(_1071_),
    .C(_1075_),
    .Y(_1079_));
 sky130_fd_sc_hd__nor2_1 _1891_ (.A(_1078_),
    .B(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__a31oi_2 _1892_ (.A1(_0924_),
    .A2(_0948_),
    .A3(_1080_),
    .B1(_1078_),
    .Y(_1081_));
 sky130_fd_sc_hd__nor2_1 _1893_ (.A(_1046_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__and2_1 _1894_ (.A(_1073_),
    .B(_1074_),
    .X(_1083_));
 sky130_fd_sc_hd__or2_1 _1895_ (.A(_1075_),
    .B(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__and3_1 _1896_ (.A(_0923_),
    .B(_0931_),
    .C(_0944_),
    .X(_1085_));
 sky130_fd_sc_hd__inv_2 _1897_ (.A(_1052_),
    .Y(_1086_));
 sky130_fd_sc_hd__o2bb2a_1 _1898_ (.A1_N(_0920_),
    .A2_N(_0938_),
    .B1(_1051_),
    .B2(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__nor2_1 _1899_ (.A(_1053_),
    .B(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__xnor2_1 _1900_ (.A(_1085_),
    .B(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__buf_2 _1901_ (.A(\MAC.a[1] ),
    .X(_1090_));
 sky130_fd_sc_hd__and3_1 _1902_ (.A(_1090_),
    .B(\MAC.a[2] ),
    .C(\MAC.b[8] ),
    .X(_1091_));
 sky130_fd_sc_hd__a21oi_1 _1903_ (.A1(\MAC.a[2] ),
    .A2(\MAC.b[8] ),
    .B1(_1090_),
    .Y(_1092_));
 sky130_fd_sc_hd__nor2_1 _1904_ (.A(_1091_),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__a31o_1 _1905_ (.A1(_0928_),
    .A2(_0939_),
    .A3(_1093_),
    .B1(_1091_),
    .X(_1094_));
 sky130_fd_sc_hd__or2b_1 _1906_ (.A(_1089_),
    .B_N(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__a21bo_1 _1907_ (.A1(_1085_),
    .A2(_1088_),
    .B1_N(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__o2bb2a_1 _1908_ (.A1_N(_0921_),
    .A2_N(_0934_),
    .B1(_1060_),
    .B2(_1061_),
    .X(_1097_));
 sky130_fd_sc_hd__nor2_1 _1909_ (.A(_1062_),
    .B(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__a22o_1 _1910_ (.A1(\MAC.a[5] ),
    .A2(_0936_),
    .B1(_0946_),
    .B2(\MAC.a[4] ),
    .X(_1099_));
 sky130_fd_sc_hd__and4_1 _1911_ (.A(\MAC.a[4] ),
    .B(\MAC.a[5] ),
    .C(\MAC.b[4] ),
    .D(_0946_),
    .X(_1100_));
 sky130_fd_sc_hd__a31o_1 _1912_ (.A1(_0914_),
    .A2(_0934_),
    .A3(_1099_),
    .B1(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__nand2_1 _1913_ (.A(_1098_),
    .B(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__xnor2_1 _1914_ (.A(_1098_),
    .B(_1101_),
    .Y(_1103_));
 sky130_fd_sc_hd__a21oi_1 _1915_ (.A1(_0923_),
    .A2(_0945_),
    .B1(_0932_),
    .Y(_1104_));
 sky130_fd_sc_hd__or2_1 _1916_ (.A(_1085_),
    .B(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__or2_1 _1917_ (.A(_1103_),
    .B(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__xnor2_1 _1918_ (.A(_0945_),
    .B(_1064_),
    .Y(_1107_));
 sky130_fd_sc_hd__a21o_1 _1919_ (.A1(_1102_),
    .A2(_1106_),
    .B1(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__or2b_1 _1920_ (.A(_1094_),
    .B_N(_1089_),
    .X(_1109_));
 sky130_fd_sc_hd__nand2_1 _1921_ (.A(_1109_),
    .B(_1095_),
    .Y(_1110_));
 sky130_fd_sc_hd__nand3_1 _1922_ (.A(_1107_),
    .B(_1102_),
    .C(_1106_),
    .Y(_1111_));
 sky130_fd_sc_hd__nand2_1 _1923_ (.A(_1108_),
    .B(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__or2_1 _1924_ (.A(_1110_),
    .B(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__xor2_1 _1925_ (.A(_1055_),
    .B(_1067_),
    .X(_1114_));
 sky130_fd_sc_hd__a21oi_1 _1926_ (.A1(_1108_),
    .A2(_1113_),
    .B1(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__and3_1 _1927_ (.A(_1114_),
    .B(_1108_),
    .C(_1113_),
    .X(_1116_));
 sky130_fd_sc_hd__nor2_1 _1928_ (.A(_1115_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__a21o_1 _1929_ (.A1(_1096_),
    .A2(_1117_),
    .B1(_1115_),
    .X(_1118_));
 sky130_fd_sc_hd__and2b_1 _1930_ (.A_N(_1084_),
    .B(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__xnor2_1 _1931_ (.A(_1084_),
    .B(_1118_),
    .Y(_1120_));
 sky130_fd_sc_hd__and3_1 _1932_ (.A(_0922_),
    .B(_0948_),
    .C(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__nand2_1 _1933_ (.A(_0924_),
    .B(_0948_),
    .Y(_1122_));
 sky130_fd_sc_hd__xnor2_1 _1934_ (.A(_1122_),
    .B(_1080_),
    .Y(_1123_));
 sky130_fd_sc_hd__o21ai_1 _1935_ (.A1(_1119_),
    .A2(_1121_),
    .B1(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__and2b_1 _1936_ (.A_N(_1100_),
    .B(_1099_),
    .X(_1125_));
 sky130_fd_sc_hd__nand2_1 _1937_ (.A(_0914_),
    .B(_0934_),
    .Y(_1126_));
 sky130_fd_sc_hd__xnor2_1 _1938_ (.A(_1125_),
    .B(_1126_),
    .Y(_1127_));
 sky130_fd_sc_hd__a22o_1 _1939_ (.A1(_0919_),
    .A2(_0936_),
    .B1(_0946_),
    .B2(_0927_),
    .X(_1128_));
 sky130_fd_sc_hd__and4_1 _1940_ (.A(_0927_),
    .B(\MAC.a[4] ),
    .C(_0936_),
    .D(_0946_),
    .X(_1129_));
 sky130_fd_sc_hd__a31o_1 _1941_ (.A1(_0912_),
    .A2(_0934_),
    .A3(_1128_),
    .B1(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__nand2_1 _1942_ (.A(_1127_),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__xor2_1 _1943_ (.A(_1127_),
    .B(_1130_),
    .X(_1132_));
 sky130_fd_sc_hd__a22o_1 _1944_ (.A1(\MAC.a[8] ),
    .A2(\MAC.b[1] ),
    .B1(\MAC.b[2] ),
    .B2(\MAC.a[7] ),
    .X(_1133_));
 sky130_fd_sc_hd__nand4_1 _1945_ (.A(\MAC.a[7] ),
    .B(\MAC.a[8] ),
    .C(_0931_),
    .D(\MAC.b[2] ),
    .Y(_1134_));
 sky130_fd_sc_hd__and3_1 _1946_ (.A(\MAC.b[0] ),
    .B(_1133_),
    .C(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__a21oi_1 _1947_ (.A1(_1133_),
    .A2(_1134_),
    .B1(\MAC.b[0] ),
    .Y(_1136_));
 sky130_fd_sc_hd__or2_1 _1948_ (.A(_1135_),
    .B(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__inv_2 _1949_ (.A(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__nand2_1 _1950_ (.A(_1132_),
    .B(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__xnor2_1 _1951_ (.A(_1103_),
    .B(_1105_),
    .Y(_1140_));
 sky130_fd_sc_hd__a21oi_1 _1952_ (.A1(_1131_),
    .A2(_1139_),
    .B1(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__and3_1 _1953_ (.A(_1140_),
    .B(_1131_),
    .C(_1139_),
    .X(_1142_));
 sky130_fd_sc_hd__or2_1 _1954_ (.A(_1141_),
    .B(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__nand2_1 _1955_ (.A(\MAC.b[8] ),
    .B(_0917_),
    .Y(_1144_));
 sky130_fd_sc_hd__a21o_1 _1956_ (.A1(\MAC.a[1] ),
    .A2(\MAC.b[8] ),
    .B1(\MAC.a[0] ),
    .X(_1145_));
 sky130_fd_sc_hd__and2_1 _1957_ (.A(_1144_),
    .B(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__nand3_1 _1958_ (.A(_0926_),
    .B(_0938_),
    .C(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__a21bo_1 _1959_ (.A1(_0930_),
    .A2(_1133_),
    .B1_N(_1134_),
    .X(_1148_));
 sky130_fd_sc_hd__nand2_1 _1960_ (.A(_0927_),
    .B(\MAC.b[7] ),
    .Y(_1149_));
 sky130_fd_sc_hd__xnor2_1 _1961_ (.A(_1093_),
    .B(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__xnor2_1 _1962_ (.A(_1148_),
    .B(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__and3_1 _1963_ (.A(_1144_),
    .B(_1147_),
    .C(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__a21oi_1 _1964_ (.A1(_1144_),
    .A2(_1147_),
    .B1(_1151_),
    .Y(_1153_));
 sky130_fd_sc_hd__or2_1 _1965_ (.A(_1152_),
    .B(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__nor2_1 _1966_ (.A(_1143_),
    .B(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__nand2_1 _1967_ (.A(_1110_),
    .B(_1112_),
    .Y(_1156_));
 sky130_fd_sc_hd__o211a_1 _1968_ (.A1(_1141_),
    .A2(_1155_),
    .B1(_1113_),
    .C1(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__and2_1 _1969_ (.A(_1148_),
    .B(_1150_),
    .X(_1158_));
 sky130_fd_sc_hd__inv_2 _1970_ (.A(_1157_),
    .Y(_1159_));
 sky130_fd_sc_hd__a211o_1 _1971_ (.A1(_1113_),
    .A2(_1156_),
    .B1(_1141_),
    .C1(_1155_),
    .X(_1160_));
 sky130_fd_sc_hd__o211a_1 _1972_ (.A1(_1158_),
    .A2(_1153_),
    .B1(_1159_),
    .C1(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__or2_1 _1973_ (.A(_1115_),
    .B(_1116_),
    .X(_1162_));
 sky130_fd_sc_hd__xnor2_1 _1974_ (.A(_1096_),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__o21a_1 _1975_ (.A1(_1157_),
    .A2(_1161_),
    .B1(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__nor3_1 _1976_ (.A(_1163_),
    .B(_1157_),
    .C(_1161_),
    .Y(_1165_));
 sky130_fd_sc_hd__nor2_1 _1977_ (.A(_1164_),
    .B(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__and3_1 _1978_ (.A(_0915_),
    .B(\MAC.b[6] ),
    .C(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__a21oi_1 _1979_ (.A1(_0922_),
    .A2(_0948_),
    .B1(_1120_),
    .Y(_1168_));
 sky130_fd_sc_hd__nor2_1 _1980_ (.A(_1121_),
    .B(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__o21ai_1 _1981_ (.A1(_1164_),
    .A2(_1167_),
    .B1(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__and4_1 _1982_ (.A(\MAC.a[2] ),
    .B(\MAC.a[3] ),
    .C(\MAC.b[4] ),
    .D(\MAC.b[5] ),
    .X(_1171_));
 sky130_fd_sc_hd__a22oi_1 _1983_ (.A1(_0927_),
    .A2(_0936_),
    .B1(_0946_),
    .B2(\MAC.a[2] ),
    .Y(_1172_));
 sky130_fd_sc_hd__and4bb_1 _1984_ (.A_N(_1171_),
    .B_N(_1172_),
    .C(_0919_),
    .D(\MAC.b[3] ),
    .X(_1173_));
 sky130_fd_sc_hd__nor2_1 _1985_ (.A(_1171_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__nand2_1 _1986_ (.A(_0912_),
    .B(_0934_),
    .Y(_1175_));
 sky130_fd_sc_hd__and2b_1 _1987_ (.A_N(_1129_),
    .B(_1128_),
    .X(_1176_));
 sky130_fd_sc_hd__xnor2_1 _1988_ (.A(_1175_),
    .B(_1176_),
    .Y(_0059_));
 sky130_fd_sc_hd__or2b_1 _1989_ (.A(_1174_),
    .B_N(_0059_),
    .X(_0060_));
 sky130_fd_sc_hd__a22oi_1 _1990_ (.A1(\MAC.a[7] ),
    .A2(_0931_),
    .B1(_0944_),
    .B2(_0914_),
    .Y(_0061_));
 sky130_fd_sc_hd__and4_1 _1991_ (.A(_0914_),
    .B(\MAC.a[7] ),
    .C(_0931_),
    .D(_0944_),
    .X(_0062_));
 sky130_fd_sc_hd__nor2_1 _1992_ (.A(_0061_),
    .B(_0062_),
    .Y(_0063_));
 sky130_fd_sc_hd__nand2_1 _1993_ (.A(_0923_),
    .B(\MAC.b[0] ),
    .Y(_0064_));
 sky130_fd_sc_hd__xnor2_1 _1994_ (.A(_0063_),
    .B(_0064_),
    .Y(_0065_));
 sky130_fd_sc_hd__xnor2_1 _1995_ (.A(_0059_),
    .B(_1174_),
    .Y(_0066_));
 sky130_fd_sc_hd__nand2_1 _1996_ (.A(_0065_),
    .B(_0066_),
    .Y(_0067_));
 sky130_fd_sc_hd__or2_1 _1997_ (.A(_1132_),
    .B(_1138_),
    .X(_0068_));
 sky130_fd_sc_hd__nand2_1 _1998_ (.A(_1139_),
    .B(_0068_),
    .Y(_0069_));
 sky130_fd_sc_hd__a21oi_2 _1999_ (.A1(_0060_),
    .A2(_0067_),
    .B1(_0069_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _2000_ (.A(_0070_),
    .Y(_0071_));
 sky130_fd_sc_hd__and3_1 _2001_ (.A(_0069_),
    .B(_0060_),
    .C(_0067_),
    .X(_0072_));
 sky130_fd_sc_hd__and3_1 _2002_ (.A(_0938_),
    .B(_0940_),
    .C(_0917_),
    .X(_0073_));
 sky130_fd_sc_hd__a31o_1 _2003_ (.A1(_0923_),
    .A2(\MAC.b[0] ),
    .A3(_0063_),
    .B1(_0062_),
    .X(_0074_));
 sky130_fd_sc_hd__nand2_1 _2004_ (.A(\MAC.a[2] ),
    .B(\MAC.b[7] ),
    .Y(_0075_));
 sky130_fd_sc_hd__xor2_1 _2005_ (.A(_1146_),
    .B(_0075_),
    .X(_0076_));
 sky130_fd_sc_hd__xnor2_1 _2006_ (.A(_0074_),
    .B(_0076_),
    .Y(_0077_));
 sky130_fd_sc_hd__nor2_1 _2007_ (.A(_0073_),
    .B(_0077_),
    .Y(_0078_));
 sky130_fd_sc_hd__and2_1 _2008_ (.A(_0073_),
    .B(_0077_),
    .X(_0079_));
 sky130_fd_sc_hd__or2_1 _2009_ (.A(_0078_),
    .B(_0079_),
    .X(_0080_));
 sky130_fd_sc_hd__or3_1 _2010_ (.A(_0070_),
    .B(_0072_),
    .C(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _2011_ (.A(_1143_),
    .B(_1154_),
    .X(_0082_));
 sky130_fd_sc_hd__a211oi_2 _2012_ (.A1(_0071_),
    .A2(_0081_),
    .B1(_1155_),
    .C1(_0082_),
    .Y(_0083_));
 sky130_fd_sc_hd__and2b_1 _2013_ (.A_N(_0076_),
    .B(_0074_),
    .X(_0084_));
 sky130_fd_sc_hd__o211a_1 _2014_ (.A1(_1155_),
    .A2(_0082_),
    .B1(_0071_),
    .C1(_0081_),
    .X(_0085_));
 sky130_fd_sc_hd__nor2_1 _2015_ (.A(_0083_),
    .B(_0085_),
    .Y(_0086_));
 sky130_fd_sc_hd__o21a_1 _2016_ (.A1(_0084_),
    .A2(_0079_),
    .B1(_0086_),
    .X(_0087_));
 sky130_fd_sc_hd__a211oi_1 _2017_ (.A1(_1159_),
    .A2(_1160_),
    .B1(_1158_),
    .C1(_1153_),
    .Y(_0088_));
 sky130_fd_sc_hd__nor2_1 _2018_ (.A(_1161_),
    .B(_0088_),
    .Y(_0089_));
 sky130_fd_sc_hd__o21a_1 _2019_ (.A1(_0083_),
    .A2(_0087_),
    .B1(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__nor3_1 _2020_ (.A(_0089_),
    .B(_0083_),
    .C(_0087_),
    .Y(_0091_));
 sky130_fd_sc_hd__nor2_1 _2021_ (.A(_0090_),
    .B(_0091_),
    .Y(_0092_));
 sky130_fd_sc_hd__and3_1 _2022_ (.A(_0913_),
    .B(_0948_),
    .C(_0092_),
    .X(_0093_));
 sky130_fd_sc_hd__a21oi_1 _2023_ (.A1(_0915_),
    .A2(_0948_),
    .B1(_1166_),
    .Y(_0094_));
 sky130_fd_sc_hd__nor2_1 _2024_ (.A(_1167_),
    .B(_0094_),
    .Y(_0095_));
 sky130_fd_sc_hd__o21ai_1 _2025_ (.A1(_0090_),
    .A2(_0093_),
    .B1(_0095_),
    .Y(_0096_));
 sky130_fd_sc_hd__buf_2 _2026_ (.A(\MAC.a[0] ),
    .X(_0097_));
 sky130_fd_sc_hd__a22oi_1 _2027_ (.A1(_1090_),
    .A2(_0938_),
    .B1(_0940_),
    .B2(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__or2_1 _2028_ (.A(_0073_),
    .B(_0098_),
    .X(_0099_));
 sky130_fd_sc_hd__and4_1 _2029_ (.A(\MAC.a[5] ),
    .B(\MAC.a[6] ),
    .C(_0931_),
    .D(_0944_),
    .X(_0100_));
 sky130_fd_sc_hd__a22oi_1 _2030_ (.A1(_0914_),
    .A2(_0931_),
    .B1(_0944_),
    .B2(_0912_),
    .Y(_0101_));
 sky130_fd_sc_hd__nor2_1 _2031_ (.A(_0100_),
    .B(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__a31o_1 _2032_ (.A1(_0921_),
    .A2(_0930_),
    .A3(_0102_),
    .B1(_0100_),
    .X(_0103_));
 sky130_fd_sc_hd__and2b_1 _2033_ (.A_N(_0099_),
    .B(_0103_),
    .X(_0104_));
 sky130_fd_sc_hd__o21ai_1 _2034_ (.A1(_0070_),
    .A2(_0072_),
    .B1(_0080_),
    .Y(_0105_));
 sky130_fd_sc_hd__o2bb2a_1 _2035_ (.A1_N(_0919_),
    .A2_N(\MAC.b[3] ),
    .B1(_1171_),
    .B2(_1172_),
    .X(_0106_));
 sky130_fd_sc_hd__and4_1 _2036_ (.A(\MAC.a[1] ),
    .B(\MAC.a[2] ),
    .C(\MAC.b[4] ),
    .D(\MAC.b[5] ),
    .X(_0107_));
 sky130_fd_sc_hd__a22oi_1 _2037_ (.A1(\MAC.a[2] ),
    .A2(_0936_),
    .B1(_0946_),
    .B2(\MAC.a[1] ),
    .Y(_0108_));
 sky130_fd_sc_hd__and4bb_1 _2038_ (.A_N(_0107_),
    .B_N(_0108_),
    .C(_0927_),
    .D(\MAC.b[3] ),
    .X(_0109_));
 sky130_fd_sc_hd__nor2_1 _2039_ (.A(_0107_),
    .B(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__or3_1 _2040_ (.A(_1173_),
    .B(_0106_),
    .C(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_1 _2041_ (.A(_0921_),
    .B(\MAC.b[0] ),
    .Y(_0112_));
 sky130_fd_sc_hd__xnor2_1 _2042_ (.A(_0102_),
    .B(_0112_),
    .Y(_0113_));
 sky130_fd_sc_hd__nor2_1 _2043_ (.A(_1173_),
    .B(_0106_),
    .Y(_0114_));
 sky130_fd_sc_hd__xnor2_1 _2044_ (.A(_0114_),
    .B(_0110_),
    .Y(_0115_));
 sky130_fd_sc_hd__nand2_1 _2045_ (.A(_0113_),
    .B(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__xnor2_1 _2046_ (.A(_0065_),
    .B(_0066_),
    .Y(_0117_));
 sky130_fd_sc_hd__a21o_1 _2047_ (.A1(_0111_),
    .A2(_0116_),
    .B1(_0117_),
    .X(_0118_));
 sky130_fd_sc_hd__xnor2_1 _2048_ (.A(_0103_),
    .B(_0099_),
    .Y(_0119_));
 sky130_fd_sc_hd__nand3_1 _2049_ (.A(_0117_),
    .B(_0111_),
    .C(_0116_),
    .Y(_0120_));
 sky130_fd_sc_hd__nand3_1 _2050_ (.A(_0118_),
    .B(_0119_),
    .C(_0120_),
    .Y(_0121_));
 sky130_fd_sc_hd__nand2_1 _2051_ (.A(_0118_),
    .B(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__a21o_1 _2052_ (.A1(_0081_),
    .A2(_0105_),
    .B1(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__nand3_1 _2053_ (.A(_0081_),
    .B(_0105_),
    .C(_0122_),
    .Y(_0124_));
 sky130_fd_sc_hd__a21boi_1 _2054_ (.A1(_0104_),
    .A2(_0123_),
    .B1_N(_0124_),
    .Y(_0125_));
 sky130_fd_sc_hd__or3_1 _2055_ (.A(_0084_),
    .B(_0079_),
    .C(_0086_),
    .X(_0126_));
 sky130_fd_sc_hd__and2b_1 _2056_ (.A_N(_0087_),
    .B(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__and2b_1 _2057_ (.A_N(_0125_),
    .B(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__xnor2_1 _2058_ (.A(_0127_),
    .B(_0125_),
    .Y(_0129_));
 sky130_fd_sc_hd__and3_1 _2059_ (.A(_0920_),
    .B(\MAC.b[6] ),
    .C(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__nand2_1 _2060_ (.A(_0913_),
    .B(\MAC.b[6] ),
    .Y(_0131_));
 sky130_fd_sc_hd__xnor2_1 _2061_ (.A(_0131_),
    .B(_0092_),
    .Y(_0132_));
 sky130_fd_sc_hd__o21a_1 _2062_ (.A1(_0128_),
    .A2(_0130_),
    .B1(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__a21oi_1 _2063_ (.A1(_0920_),
    .A2(\MAC.b[6] ),
    .B1(_0129_),
    .Y(_0134_));
 sky130_fd_sc_hd__or2_1 _2064_ (.A(_0130_),
    .B(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__and3_1 _2065_ (.A(_0104_),
    .B(_0124_),
    .C(_0123_),
    .X(_0136_));
 sky130_fd_sc_hd__a21oi_1 _2066_ (.A1(_0124_),
    .A2(_0123_),
    .B1(_0104_),
    .Y(_0137_));
 sky130_fd_sc_hd__or2_1 _2067_ (.A(_0136_),
    .B(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__a21o_1 _2068_ (.A1(_0118_),
    .A2(_0120_),
    .B1(_0119_),
    .X(_0139_));
 sky130_fd_sc_hd__o2bb2a_1 _2069_ (.A1_N(_0927_),
    .A2_N(_0934_),
    .B1(_0107_),
    .B2(_0108_),
    .X(_0140_));
 sky130_fd_sc_hd__and4_1 _2070_ (.A(\MAC.a[0] ),
    .B(\MAC.a[1] ),
    .C(_0936_),
    .D(_0946_),
    .X(_0141_));
 sky130_fd_sc_hd__a22oi_1 _2071_ (.A1(\MAC.a[1] ),
    .A2(_0936_),
    .B1(_0946_),
    .B2(\MAC.a[0] ),
    .Y(_0142_));
 sky130_fd_sc_hd__and4bb_1 _2072_ (.A_N(_0141_),
    .B_N(_0142_),
    .C(\MAC.a[2] ),
    .D(\MAC.b[3] ),
    .X(_0143_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(_0141_),
    .B(_0143_),
    .Y(_0144_));
 sky130_fd_sc_hd__or3_1 _2074_ (.A(_0109_),
    .B(_0140_),
    .C(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__a22oi_1 _2075_ (.A1(_0912_),
    .A2(_0931_),
    .B1(_0944_),
    .B2(_0919_),
    .Y(_0146_));
 sky130_fd_sc_hd__and4_1 _2076_ (.A(_0919_),
    .B(_0912_),
    .C(_0931_),
    .D(_0944_),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_1 _2077_ (.A(_0146_),
    .B(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__nand2_1 _2078_ (.A(_0914_),
    .B(\MAC.b[0] ),
    .Y(_0149_));
 sky130_fd_sc_hd__xnor2_1 _2079_ (.A(_0148_),
    .B(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__nor2_1 _2080_ (.A(_0109_),
    .B(_0140_),
    .Y(_0151_));
 sky130_fd_sc_hd__xnor2_1 _2081_ (.A(_0151_),
    .B(_0144_),
    .Y(_0152_));
 sky130_fd_sc_hd__nand2_1 _2082_ (.A(_0150_),
    .B(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__xnor2_1 _2083_ (.A(_0113_),
    .B(_0115_),
    .Y(_0154_));
 sky130_fd_sc_hd__a21oi_1 _2084_ (.A1(_0145_),
    .A2(_0153_),
    .B1(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__nand2_1 _2085_ (.A(_0097_),
    .B(_0938_),
    .Y(_0156_));
 sky130_fd_sc_hd__o21ba_1 _2086_ (.A1(_0146_),
    .A2(_0149_),
    .B1_N(_0147_),
    .X(_0157_));
 sky130_fd_sc_hd__xnor2_1 _2087_ (.A(_0156_),
    .B(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__and3_1 _2088_ (.A(_0154_),
    .B(_0145_),
    .C(_0153_),
    .X(_0159_));
 sky130_fd_sc_hd__or3_1 _2089_ (.A(_0155_),
    .B(_0158_),
    .C(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__or2b_1 _2090_ (.A(_0155_),
    .B_N(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__nor2_1 _2091_ (.A(_0156_),
    .B(_0157_),
    .Y(_0162_));
 sky130_fd_sc_hd__nand2_1 _2092_ (.A(_0121_),
    .B(_0139_),
    .Y(_0163_));
 sky130_fd_sc_hd__xnor2_1 _2093_ (.A(_0163_),
    .B(_0161_),
    .Y(_0164_));
 sky130_fd_sc_hd__and2_1 _2094_ (.A(_0162_),
    .B(_0164_),
    .X(_0165_));
 sky130_fd_sc_hd__a31oi_2 _2095_ (.A1(_0121_),
    .A2(_0139_),
    .A3(_0161_),
    .B1(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__xnor2_1 _2096_ (.A(_0138_),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__nand2_1 _2097_ (.A(_0928_),
    .B(\MAC.b[6] ),
    .Y(_0168_));
 sky130_fd_sc_hd__or2_1 _2098_ (.A(_0167_),
    .B(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__o21ai_1 _2099_ (.A1(_0138_),
    .A2(_0166_),
    .B1(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__and2b_1 _2100_ (.A_N(_0135_),
    .B(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__nand2_1 _2101_ (.A(_0167_),
    .B(_0168_),
    .Y(_0172_));
 sky130_fd_sc_hd__and2_1 _2102_ (.A(_0169_),
    .B(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__nor2_1 _2103_ (.A(_0162_),
    .B(_0164_),
    .Y(_0174_));
 sky130_fd_sc_hd__o2bb2a_1 _2104_ (.A1_N(_0926_),
    .A2_N(_0934_),
    .B1(_0141_),
    .B2(_0142_),
    .X(_0175_));
 sky130_fd_sc_hd__nor2_1 _2105_ (.A(_0143_),
    .B(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__and3_1 _2106_ (.A(_0935_),
    .B(_0937_),
    .C(_0917_),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _2107_ (.A(_0176_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__xnor2_1 _2108_ (.A(_0176_),
    .B(_0177_),
    .Y(_0179_));
 sky130_fd_sc_hd__nand2_1 _2109_ (.A(_0912_),
    .B(_0930_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_1 _2110_ (.A(_0919_),
    .B(_0932_),
    .Y(_0181_));
 sky130_fd_sc_hd__nand2_1 _2111_ (.A(_0927_),
    .B(_0944_),
    .Y(_0182_));
 sky130_fd_sc_hd__and4_1 _2112_ (.A(_0927_),
    .B(_0919_),
    .C(_0931_),
    .D(_0944_),
    .X(_0183_));
 sky130_fd_sc_hd__a21o_1 _2113_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__xor2_1 _2114_ (.A(_0180_),
    .B(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__or2b_1 _2115_ (.A(_0179_),
    .B_N(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__or2_1 _2116_ (.A(_0150_),
    .B(_0152_),
    .X(_0187_));
 sky130_fd_sc_hd__nand2_1 _2117_ (.A(_0153_),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__a21oi_1 _2118_ (.A1(_0178_),
    .A2(_0186_),
    .B1(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__o21ba_1 _2119_ (.A1(_0180_),
    .A2(_0184_),
    .B1_N(_0183_),
    .X(_0190_));
 sky130_fd_sc_hd__and3_1 _2120_ (.A(_0188_),
    .B(_0178_),
    .C(_0186_),
    .X(_0191_));
 sky130_fd_sc_hd__nor2_1 _2121_ (.A(_0189_),
    .B(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__and2b_1 _2122_ (.A_N(_0190_),
    .B(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__o21ai_1 _2123_ (.A1(_0155_),
    .A2(_0159_),
    .B1(_0158_),
    .Y(_0194_));
 sky130_fd_sc_hd__o211a_1 _2124_ (.A1(_0189_),
    .A2(_0193_),
    .B1(_0160_),
    .C1(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__or3b_1 _2125_ (.A(_0165_),
    .B(_0174_),
    .C_N(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__nand2_1 _2126_ (.A(_0926_),
    .B(\MAC.b[6] ),
    .Y(_0197_));
 sky130_fd_sc_hd__or2_1 _2127_ (.A(_0165_),
    .B(_0174_),
    .X(_0198_));
 sky130_fd_sc_hd__xor2_1 _2128_ (.A(_0198_),
    .B(_0195_),
    .X(_0199_));
 sky130_fd_sc_hd__or2_1 _2129_ (.A(_0197_),
    .B(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__nand2_1 _2130_ (.A(_0196_),
    .B(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__nand2_1 _2131_ (.A(_0173_),
    .B(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__xnor2_1 _2132_ (.A(_0173_),
    .B(_0201_),
    .Y(_0203_));
 sky130_fd_sc_hd__xnor2_1 _2133_ (.A(_0179_),
    .B(_0185_),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_2 _2134_ (.A(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__a22o_1 _2135_ (.A1(_0928_),
    .A2(_0932_),
    .B1(_0945_),
    .B2(_0926_),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_1 _2136_ (.A(\MAC.a[2] ),
    .B(_0932_),
    .Y(_0207_));
 sky130_fd_sc_hd__or2_1 _2137_ (.A(_0182_),
    .B(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__nand2_1 _2138_ (.A(_0206_),
    .B(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__nand2_1 _2139_ (.A(_0919_),
    .B(_0930_),
    .Y(_0210_));
 sky130_fd_sc_hd__xor2_1 _2140_ (.A(_0209_),
    .B(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__a22o_1 _2141_ (.A1(_1090_),
    .A2(_0935_),
    .B1(_0937_),
    .B2(_0097_),
    .X(_0212_));
 sky130_fd_sc_hd__nand3b_1 _2142_ (.A_N(_0177_),
    .B(_0211_),
    .C(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__xor2_1 _2143_ (.A(_0204_),
    .B(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__o21ai_1 _2144_ (.A1(_0209_),
    .A2(_0210_),
    .B1(_0208_),
    .Y(_0215_));
 sky130_fd_sc_hd__and2b_1 _2145_ (.A_N(_0214_),
    .B(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__o21ba_1 _2146_ (.A1(_0205_),
    .A2(_0213_),
    .B1_N(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__xnor2_1 _2147_ (.A(_0190_),
    .B(_0192_),
    .Y(_0218_));
 sky130_fd_sc_hd__or2b_1 _2148_ (.A(_0217_),
    .B_N(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__a211oi_1 _2149_ (.A1(_0160_),
    .A2(_0194_),
    .B1(_0189_),
    .C1(_0193_),
    .Y(_0220_));
 sky130_fd_sc_hd__or3_1 _2150_ (.A(_0195_),
    .B(_0219_),
    .C(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__and2_1 _2151_ (.A(_1090_),
    .B(\MAC.b[6] ),
    .X(_0222_));
 sky130_fd_sc_hd__o21ai_1 _2152_ (.A1(_0195_),
    .A2(_0220_),
    .B1(_0219_),
    .Y(_0223_));
 sky130_fd_sc_hd__nand3_1 _2153_ (.A(_0221_),
    .B(_0222_),
    .C(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__a21o_1 _2154_ (.A1(_0221_),
    .A2(_0223_),
    .B1(_0222_),
    .X(_0225_));
 sky130_fd_sc_hd__xnor2_1 _2155_ (.A(_0218_),
    .B(_0217_),
    .Y(_0226_));
 sky130_fd_sc_hd__a21o_1 _2156_ (.A1(_0097_),
    .A2(\MAC.b[6] ),
    .B1(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__xnor2_1 _2157_ (.A(_0215_),
    .B(_0214_),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_1 _2158_ (.A(_1090_),
    .B(_0945_),
    .Y(_0229_));
 sky130_fd_sc_hd__and4_1 _2159_ (.A(_1090_),
    .B(_0926_),
    .C(_0932_),
    .D(_0945_),
    .X(_0230_));
 sky130_fd_sc_hd__a21oi_1 _2160_ (.A1(_0207_),
    .A2(_0229_),
    .B1(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__nand2_1 _2161_ (.A(_0928_),
    .B(_0930_),
    .Y(_0232_));
 sky130_fd_sc_hd__xnor2_1 _2162_ (.A(_0231_),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__and3_1 _2163_ (.A(_0097_),
    .B(_0935_),
    .C(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__and4b_1 _2164_ (.A_N(_0231_),
    .B(_0917_),
    .C(_0932_),
    .D(_0930_),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_1 _2165_ (.A1(_1090_),
    .A2(_0932_),
    .B1(_0945_),
    .B2(_0097_),
    .X(_0236_));
 sky130_fd_sc_hd__and4_1 _2166_ (.A(_0097_),
    .B(_1090_),
    .C(_0932_),
    .D(_0945_),
    .X(_0237_));
 sky130_fd_sc_hd__a31o_1 _2167_ (.A1(_0926_),
    .A2(_0930_),
    .A3(_0236_),
    .B1(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__or3_1 _2168_ (.A(_0234_),
    .B(_0235_),
    .C(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__and2_1 _2169_ (.A(_0235_),
    .B(_0238_),
    .X(_0240_));
 sky130_fd_sc_hd__a211o_1 _2170_ (.A1(_0097_),
    .A2(_0935_),
    .B1(_0233_),
    .C1(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__a31o_1 _2171_ (.A1(_0928_),
    .A2(_0930_),
    .A3(_0231_),
    .B1(_0230_),
    .X(_0242_));
 sky130_fd_sc_hd__or2b_1 _2172_ (.A(_0177_),
    .B_N(_0212_),
    .X(_0243_));
 sky130_fd_sc_hd__xnor2_1 _2173_ (.A(_0211_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__a32o_1 _2174_ (.A1(_0228_),
    .A2(_0239_),
    .A3(_0241_),
    .B1(_0242_),
    .B2(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__or2_1 _2175_ (.A(_0244_),
    .B(_0242_),
    .X(_0246_));
 sky130_fd_sc_hd__a22o_1 _2176_ (.A1(_0234_),
    .A2(_0240_),
    .B1(_0246_),
    .B2(_0228_),
    .X(_0247_));
 sky130_fd_sc_hd__a32o_1 _2177_ (.A1(_0097_),
    .A2(\MAC.b[6] ),
    .A3(_0226_),
    .B1(_0245_),
    .B2(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__nand4_1 _2178_ (.A(_0225_),
    .B(_0227_),
    .C(_0248_),
    .D(_0224_),
    .Y(_0249_));
 sky130_fd_sc_hd__nand2_1 _2179_ (.A(_0197_),
    .B(_0199_),
    .Y(_0250_));
 sky130_fd_sc_hd__o2bb2a_1 _2180_ (.A1_N(_0200_),
    .A2_N(_0250_),
    .B1(_0221_),
    .B2(_0249_),
    .X(_0251_));
 sky130_fd_sc_hd__a31o_1 _2181_ (.A1(_0221_),
    .A2(_0224_),
    .A3(_0249_),
    .B1(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__or2_1 _2182_ (.A(_0203_),
    .B(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__xor2_1 _2183_ (.A(_0135_),
    .B(_0170_),
    .X(_0254_));
 sky130_fd_sc_hd__a21oi_1 _2184_ (.A1(_0202_),
    .A2(_0253_),
    .B1(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__nor3_1 _2185_ (.A(_0132_),
    .B(_0128_),
    .C(_0130_),
    .Y(_0256_));
 sky130_fd_sc_hd__nor2_1 _2186_ (.A(_0133_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__o21a_1 _2187_ (.A1(_0171_),
    .A2(_0255_),
    .B1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__or3_1 _2188_ (.A(_0095_),
    .B(_0090_),
    .C(_0093_),
    .X(_0259_));
 sky130_fd_sc_hd__and2_1 _2189_ (.A(_0096_),
    .B(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__o21ai_1 _2190_ (.A1(_0133_),
    .A2(_0258_),
    .B1(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__or3_1 _2191_ (.A(_1169_),
    .B(_1164_),
    .C(_1167_),
    .X(_0262_));
 sky130_fd_sc_hd__nand2_1 _2192_ (.A(_1170_),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__a21o_1 _2193_ (.A1(_0096_),
    .A2(_0261_),
    .B1(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__or3_1 _2194_ (.A(_1123_),
    .B(_1119_),
    .C(_1121_),
    .X(_0265_));
 sky130_fd_sc_hd__nand2_1 _2195_ (.A(_1124_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__a21o_1 _2196_ (.A1(_1170_),
    .A2(_0264_),
    .B1(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__xnor2_1 _2197_ (.A(_1046_),
    .B(_1081_),
    .Y(_0268_));
 sky130_fd_sc_hd__a21oi_1 _2198_ (.A1(_1124_),
    .A2(_0267_),
    .B1(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__nor3_1 _2199_ (.A(_1043_),
    .B(_1038_),
    .C(_1041_),
    .Y(_0270_));
 sky130_fd_sc_hd__nor2_1 _2200_ (.A(_1044_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__o21a_1 _2201_ (.A1(_1082_),
    .A2(_0269_),
    .B1(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_1 _2202_ (.A(_1044_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__o21ai_1 _2203_ (.A1(_1013_),
    .A2(_0273_),
    .B1(_1011_),
    .Y(_0274_));
 sky130_fd_sc_hd__and3b_1 _2204_ (.A_N(_0957_),
    .B(_0965_),
    .C(_0956_),
    .X(_0275_));
 sky130_fd_sc_hd__or3b_1 _2205_ (.A(_0981_),
    .B(_0274_),
    .C_N(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__buf_2 _2206_ (.A(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__inv_2 _2207_ (.A(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand2_1 _2208_ (.A(_0203_),
    .B(_0252_),
    .Y(_0279_));
 sky130_fd_sc_hd__nand2_1 _2209_ (.A(_0253_),
    .B(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__or4_1 _2210_ (.A(_0945_),
    .B(_0935_),
    .C(_0937_),
    .D(_0947_),
    .X(_0281_));
 sky130_fd_sc_hd__or4_1 _2211_ (.A(\MAC.b[14] ),
    .B(\MAC.b[13] ),
    .C(_0930_),
    .D(_0932_),
    .X(_0282_));
 sky130_fd_sc_hd__or4_1 _2212_ (.A(\MAC.b[10] ),
    .B(\MAC.b[9] ),
    .C(\MAC.b[12] ),
    .D(\MAC.b[11] ),
    .X(_0283_));
 sky130_fd_sc_hd__or4_1 _2213_ (.A(_0948_),
    .B(_0939_),
    .C(_0941_),
    .D(\MAC.b[15] ),
    .X(_0284_));
 sky130_fd_sc_hd__or3_1 _2214_ (.A(_0282_),
    .B(_0283_),
    .C(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__or4_1 _2215_ (.A(\MAC.a[12] ),
    .B(\MAC.a[11] ),
    .C(\MAC.a[14] ),
    .D(\MAC.a[13] ),
    .X(_0286_));
 sky130_fd_sc_hd__or4_1 _2216_ (.A(\MAC.a[10] ),
    .B(\MAC.a[9] ),
    .C(_0920_),
    .D(_0913_),
    .X(_0287_));
 sky130_fd_sc_hd__or4_1 _2217_ (.A(_0097_),
    .B(_1090_),
    .C(_0926_),
    .D(_0928_),
    .X(_0288_));
 sky130_fd_sc_hd__or4_1 _2218_ (.A(_0915_),
    .B(_0922_),
    .C(_0924_),
    .D(\MAC.a[15] ),
    .X(_0289_));
 sky130_fd_sc_hd__or4_1 _2219_ (.A(_0286_),
    .B(_0287_),
    .C(_0288_),
    .D(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__o21a_2 _2220_ (.A1(_0281_),
    .A2(_0285_),
    .B1(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__inv_2 _2221_ (.A(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__and3_1 _2222_ (.A(_0254_),
    .B(_0202_),
    .C(_0253_),
    .X(_0293_));
 sky130_fd_sc_hd__nor2_1 _2223_ (.A(_0255_),
    .B(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__nor2_1 _2224_ (.A(_0278_),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__a211o_1 _2225_ (.A1(_0278_),
    .A2(_0280_),
    .B1(_0292_),
    .C1(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__inv_2 _2226_ (.A(_0891_),
    .Y(_0297_));
 sky130_fd_sc_hd__or3_1 _2227_ (.A(_0881_),
    .B(_0887_),
    .C(_0904_),
    .X(_0298_));
 sky130_fd_sc_hd__nor2_1 _2228_ (.A(_0297_),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__xnor2_1 _2229_ (.A(_0897_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2_1 _2230_ (.A(_0895_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__or2_1 _2231_ (.A(_0878_),
    .B(_0893_),
    .X(_0302_));
 sky130_fd_sc_hd__buf_2 _2232_ (.A(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__nand2_1 _2233_ (.A(_0301_),
    .B(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__a21oi_1 _2234_ (.A1(_0952_),
    .A2(_0296_),
    .B1(_0304_),
    .Y(\MAC.mul.c_mul1[0] ));
 sky130_fd_sc_hd__nor3_1 _2235_ (.A(_0257_),
    .B(_0171_),
    .C(_0255_),
    .Y(_0305_));
 sky130_fd_sc_hd__nor2_1 _2236_ (.A(_0258_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__mux2_1 _2237_ (.A0(_0294_),
    .A1(_0306_),
    .S(_0277_),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_1 _2238_ (.A(_0301_),
    .B(_0952_),
    .Y(_0308_));
 sky130_fd_sc_hd__buf_2 _2239_ (.A(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__a21o_1 _2240_ (.A1(_0291_),
    .A2(_0307_),
    .B1(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__and2_1 _2241_ (.A(_0303_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__clkbuf_1 _2242_ (.A(_0311_),
    .X(\MAC.mul.c_mul1[1] ));
 sky130_fd_sc_hd__or3_1 _2243_ (.A(_0260_),
    .B(_0133_),
    .C(_0258_),
    .X(_0312_));
 sky130_fd_sc_hd__and2_1 _2244_ (.A(_0261_),
    .B(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2245_ (.A0(_0306_),
    .A1(_0313_),
    .S(_0277_),
    .X(_0314_));
 sky130_fd_sc_hd__a21o_1 _2246_ (.A1(_0291_),
    .A2(_0314_),
    .B1(_0309_),
    .X(_0315_));
 sky130_fd_sc_hd__and2_1 _2247_ (.A(_0303_),
    .B(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_1 _2248_ (.A(_0316_),
    .X(\MAC.mul.c_mul1[2] ));
 sky130_fd_sc_hd__nand3_1 _2249_ (.A(_0263_),
    .B(_0096_),
    .C(_0261_),
    .Y(_0317_));
 sky130_fd_sc_hd__and2_1 _2250_ (.A(_0264_),
    .B(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2251_ (.A0(_0313_),
    .A1(_0318_),
    .S(_0277_),
    .X(_0319_));
 sky130_fd_sc_hd__a21o_1 _2252_ (.A1(_0291_),
    .A2(_0319_),
    .B1(_0309_),
    .X(_0320_));
 sky130_fd_sc_hd__and2_1 _2253_ (.A(_0303_),
    .B(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _2254_ (.A(_0321_),
    .X(\MAC.mul.c_mul1[3] ));
 sky130_fd_sc_hd__nand3_1 _2255_ (.A(_0266_),
    .B(_1170_),
    .C(_0264_),
    .Y(_0322_));
 sky130_fd_sc_hd__and2_1 _2256_ (.A(_0267_),
    .B(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _2257_ (.A0(_0318_),
    .A1(_0323_),
    .S(_0277_),
    .X(_0324_));
 sky130_fd_sc_hd__a21o_1 _2258_ (.A1(_0291_),
    .A2(_0324_),
    .B1(_0309_),
    .X(_0325_));
 sky130_fd_sc_hd__and2_1 _2259_ (.A(_0303_),
    .B(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _2260_ (.A(_0326_),
    .X(\MAC.mul.c_mul1[4] ));
 sky130_fd_sc_hd__buf_2 _2261_ (.A(_0277_),
    .X(_0327_));
 sky130_fd_sc_hd__and3_1 _2262_ (.A(_0268_),
    .B(_1124_),
    .C(_0267_),
    .X(_0328_));
 sky130_fd_sc_hd__or2_1 _2263_ (.A(_0269_),
    .B(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _2264_ (.A(_0327_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__o211a_1 _2265_ (.A1(_0327_),
    .A2(_0323_),
    .B1(_0330_),
    .C1(_0291_),
    .X(_0331_));
 sky130_fd_sc_hd__o21a_1 _2266_ (.A1(_0309_),
    .A2(_0331_),
    .B1(_0303_),
    .X(\MAC.mul.c_mul1[5] ));
 sky130_fd_sc_hd__nor3_1 _2267_ (.A(_1082_),
    .B(_0269_),
    .C(_0271_),
    .Y(_0332_));
 sky130_fd_sc_hd__or2_1 _2268_ (.A(_0272_),
    .B(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _2269_ (.A0(_0329_),
    .A1(_0333_),
    .S(_0327_),
    .X(_0334_));
 sky130_fd_sc_hd__nor2_1 _2270_ (.A(_0292_),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__o21a_1 _2271_ (.A1(_0309_),
    .A2(_0335_),
    .B1(_0303_),
    .X(\MAC.mul.c_mul1[6] ));
 sky130_fd_sc_hd__xnor2_1 _2272_ (.A(_1013_),
    .B(_0273_),
    .Y(_0336_));
 sky130_fd_sc_hd__mux2_1 _2273_ (.A0(_0333_),
    .A1(_0336_),
    .S(_0327_),
    .X(_0337_));
 sky130_fd_sc_hd__nor2_1 _2274_ (.A(_0292_),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__o21a_1 _2275_ (.A1(_0309_),
    .A2(_0338_),
    .B1(_0303_),
    .X(\MAC.mul.c_mul1[7] ));
 sky130_fd_sc_hd__or2_1 _2276_ (.A(_0327_),
    .B(_0336_),
    .X(_0339_));
 sky130_fd_sc_hd__a41o_1 _2277_ (.A1(_0922_),
    .A2(_0924_),
    .A3(_0939_),
    .A4(_0941_),
    .B1(_0275_),
    .X(_0340_));
 sky130_fd_sc_hd__xnor2_1 _2278_ (.A(_0981_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__xnor2_1 _2279_ (.A(_0274_),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _2280_ (.A(_0327_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__a21oi_1 _2281_ (.A1(_0339_),
    .A2(_0343_),
    .B1(_0292_),
    .Y(_0344_));
 sky130_fd_sc_hd__o21a_1 _2282_ (.A1(_0309_),
    .A2(_0344_),
    .B1(_0303_),
    .X(\MAC.mul.c_mul1[8] ));
 sky130_fd_sc_hd__and2_1 _2283_ (.A(_0885_),
    .B(_0902_),
    .X(_0345_));
 sky130_fd_sc_hd__or2_1 _2284_ (.A(_0345_),
    .B(_0327_),
    .X(_0346_));
 sky130_fd_sc_hd__nand2_1 _2285_ (.A(_0345_),
    .B(_0327_),
    .Y(_0347_));
 sky130_fd_sc_hd__a21o_1 _2286_ (.A1(_0346_),
    .A2(_0347_),
    .B1(_0292_),
    .X(_0348_));
 sky130_fd_sc_hd__a21oi_1 _2287_ (.A1(_0952_),
    .A2(_0348_),
    .B1(_0304_),
    .Y(\MAC.mul.c_mul1[9] ));
 sky130_fd_sc_hd__o21a_1 _2288_ (.A1(_0345_),
    .A2(_0327_),
    .B1(_0909_),
    .X(_0349_));
 sky130_fd_sc_hd__or3_1 _2289_ (.A(_0345_),
    .B(_0909_),
    .C(_0327_),
    .X(_0350_));
 sky130_fd_sc_hd__and3b_1 _2290_ (.A_N(_0349_),
    .B(_0350_),
    .C(_0291_),
    .X(_0351_));
 sky130_fd_sc_hd__o21a_1 _2291_ (.A1(_0309_),
    .A2(_0351_),
    .B1(_0303_),
    .X(\MAC.mul.c_mul1[10] ));
 sky130_fd_sc_hd__or3b_2 _2292_ (.A(_0907_),
    .B(_0910_),
    .C_N(_0277_),
    .X(_0352_));
 sky130_fd_sc_hd__o21ai_1 _2293_ (.A1(_0910_),
    .A2(_0278_),
    .B1(_0907_),
    .Y(_0353_));
 sky130_fd_sc_hd__a31o_1 _2294_ (.A1(_0291_),
    .A2(_0352_),
    .A3(_0353_),
    .B1(_0308_),
    .X(_0354_));
 sky130_fd_sc_hd__and2_1 _2295_ (.A(_0302_),
    .B(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _2296_ (.A(_0355_),
    .X(\MAC.mul.c_mul1[11] ));
 sky130_fd_sc_hd__or2b_1 _2297_ (.A(_0904_),
    .B_N(_0906_),
    .X(_0356_));
 sky130_fd_sc_hd__a21oi_1 _2298_ (.A1(_0356_),
    .A2(_0352_),
    .B1(_0901_),
    .Y(_0357_));
 sky130_fd_sc_hd__a31o_1 _2299_ (.A1(_0901_),
    .A2(_0356_),
    .A3(_0352_),
    .B1(_0292_),
    .X(_0358_));
 sky130_fd_sc_hd__o21bai_1 _2300_ (.A1(_0357_),
    .A2(_0358_),
    .B1_N(_0308_),
    .Y(_0359_));
 sky130_fd_sc_hd__and2_1 _2301_ (.A(_0302_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _2302_ (.A(_0360_),
    .X(\MAC.mul.c_mul1[12] ));
 sky130_fd_sc_hd__a21o_1 _2303_ (.A1(_0298_),
    .A2(_0899_),
    .B1(_0299_),
    .X(_0361_));
 sky130_fd_sc_hd__or3_1 _2304_ (.A(_0901_),
    .B(_0352_),
    .C(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__o21ai_1 _2305_ (.A1(_0901_),
    .A2(_0352_),
    .B1(_0361_),
    .Y(_0363_));
 sky130_fd_sc_hd__a31o_1 _2306_ (.A1(_0291_),
    .A2(_0362_),
    .A3(_0363_),
    .B1(_0308_),
    .X(_0364_));
 sky130_fd_sc_hd__and2_1 _2307_ (.A(_0302_),
    .B(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _2308_ (.A(_0365_),
    .X(\MAC.mul.c_mul1[13] ));
 sky130_fd_sc_hd__xor2_1 _2309_ (.A(_0300_),
    .B(_0362_),
    .X(_0366_));
 sky130_fd_sc_hd__a21o_1 _2310_ (.A1(_0291_),
    .A2(_0366_),
    .B1(_0309_),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _2311_ (.A(_0302_),
    .B(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _2312_ (.A(_0368_),
    .X(\MAC.mul.c_mul1[14] ));
 sky130_fd_sc_hd__nor2_1 _2313_ (.A(\MAC.a[15] ),
    .B(\MAC.b[15] ),
    .Y(_0369_));
 sky130_fd_sc_hd__and2_1 _2314_ (.A(\MAC.a[15] ),
    .B(\MAC.b[15] ),
    .X(_0370_));
 sky130_fd_sc_hd__or3_1 _2315_ (.A(_0292_),
    .B(_0369_),
    .C(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__a21oi_1 _2316_ (.A1(_0952_),
    .A2(_0371_),
    .B1(_0304_),
    .Y(\MAC.mul.c_mul1[15] ));
 sky130_fd_sc_hd__mux2_1 _2317_ (.A0(\MAC.add.b1[8] ),
    .A1(\MAC.add.b1[0] ),
    .S(\wrap2.state[0] ),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_1 _2318_ (.A(_0372_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2319_ (.A0(\MAC.add.b1[9] ),
    .A1(\MAC.add.b1[1] ),
    .S(\wrap2.state[0] ),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _2320_ (.A(_0373_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2321_ (.A0(\MAC.add.b1[10] ),
    .A1(\MAC.add.b1[2] ),
    .S(\wrap2.state[0] ),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _2322_ (.A(_0374_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2323_ (.A0(\MAC.add.b1[11] ),
    .A1(\MAC.add.b1[3] ),
    .S(\wrap2.state[0] ),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _2324_ (.A(_0375_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2325_ (.A0(\MAC.add.b1[12] ),
    .A1(\MAC.add.b1[4] ),
    .S(\wrap2.state[0] ),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _2326_ (.A(_0376_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2327_ (.A0(\MAC.add.b1[13] ),
    .A1(\MAC.add.b1[5] ),
    .S(\wrap2.state[0] ),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _2328_ (.A(_0377_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2329_ (.A0(\MAC.add.b1[14] ),
    .A1(\MAC.add.b1[6] ),
    .S(\wrap2.state[0] ),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _2330_ (.A(_0378_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2331_ (.A0(\MAC.add.b1[15] ),
    .A1(\MAC.add.b1[7] ),
    .S(\wrap2.state[0] ),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_1 _2332_ (.A(_0379_),
    .X(_0041_));
 sky130_fd_sc_hd__or3_1 _2333_ (.A(_0657_),
    .B(_0538_),
    .C(_0837_),
    .X(_0380_));
 sky130_fd_sc_hd__inv_2 _2334_ (.A(\MAC.add.a1[4] ),
    .Y(_0381_));
 sky130_fd_sc_hd__inv_2 _2335_ (.A(\MAC.add.a1[5] ),
    .Y(_0382_));
 sky130_fd_sc_hd__a22o_1 _2336_ (.A1(_0381_),
    .A2(\MAC.add.b1[4] ),
    .B1(_0382_),
    .B2(\MAC.add.b1[5] ),
    .X(_0383_));
 sky130_fd_sc_hd__inv_2 _2337_ (.A(\MAC.add.a1[3] ),
    .Y(_0384_));
 sky130_fd_sc_hd__inv_2 _2338_ (.A(\MAC.add.a1[2] ),
    .Y(_0385_));
 sky130_fd_sc_hd__a2bb2o_1 _2339_ (.A1_N(_0384_),
    .A2_N(\MAC.add.b1[3] ),
    .B1(_0385_),
    .B2(\MAC.add.b1[2] ),
    .X(_0386_));
 sky130_fd_sc_hd__a221o_1 _2340_ (.A1(_0551_),
    .A2(\MAC.add.b1[0] ),
    .B1(_0576_),
    .B2(\MAC.add.b1[1] ),
    .C1(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__inv_2 _2341_ (.A(\MAC.add.a1[6] ),
    .Y(_0388_));
 sky130_fd_sc_hd__and2_1 _2342_ (.A(_0388_),
    .B(\MAC.add.b1[6] ),
    .X(_0389_));
 sky130_fd_sc_hd__and2_1 _2343_ (.A(_0384_),
    .B(\MAC.add.b1[3] ),
    .X(_0390_));
 sky130_fd_sc_hd__a21o_1 _2344_ (.A1(\MAC.add.a1[1] ),
    .A2(_0577_),
    .B1(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__nor2_1 _2345_ (.A(_0382_),
    .B(\MAC.add.b1[5] ),
    .Y(_0392_));
 sky130_fd_sc_hd__or2_1 _2346_ (.A(_0385_),
    .B(\MAC.add.b1[2] ),
    .X(_0393_));
 sky130_fd_sc_hd__inv_2 _2347_ (.A(\MAC.add.a1[7] ),
    .Y(_0394_));
 sky130_fd_sc_hd__and2_1 _2348_ (.A(_0394_),
    .B(\MAC.add.b1[7] ),
    .X(_0395_));
 sky130_fd_sc_hd__a21oi_1 _2349_ (.A1(\MAC.add.a1[0] ),
    .A2(_0552_),
    .B1(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__o211a_1 _2350_ (.A1(_0381_),
    .A2(\MAC.add.b1[4] ),
    .B1(_0393_),
    .C1(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__or4b_1 _2351_ (.A(_0389_),
    .B(_0391_),
    .C(_0392_),
    .D_N(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__o22a_1 _2352_ (.A1(_0388_),
    .A2(\MAC.add.b1[6] ),
    .B1(_0394_),
    .B2(\MAC.add.b1[7] ),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_1 _2353_ (.A(_0567_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__inv_2 _2354_ (.A(\MAC.add.a1[8] ),
    .Y(_0401_));
 sky130_fd_sc_hd__or3_1 _2355_ (.A(_0576_),
    .B(\MAC.add.b1[1] ),
    .C(_0386_),
    .X(_0402_));
 sky130_fd_sc_hd__a31o_1 _2356_ (.A1(_0387_),
    .A2(_0402_),
    .A3(_0393_),
    .B1(_0390_),
    .X(_0403_));
 sky130_fd_sc_hd__o221a_1 _2357_ (.A1(_0384_),
    .A2(\MAC.add.b1[3] ),
    .B1(_0381_),
    .B2(\MAC.add.b1[4] ),
    .C1(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__o21ba_1 _2358_ (.A1(_0383_),
    .A2(_0404_),
    .B1_N(_0392_),
    .X(_0405_));
 sky130_fd_sc_hd__or2_1 _2359_ (.A(_0389_),
    .B(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__a221o_1 _2360_ (.A1(\MAC.add.b1[8] ),
    .A2(_0401_),
    .B1(_0399_),
    .B2(_0406_),
    .C1(_0395_),
    .X(_0407_));
 sky130_fd_sc_hd__o21ai_1 _2361_ (.A1(\MAC.add.b1[8] ),
    .A2(_0401_),
    .B1(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__o41a_1 _2362_ (.A1(_0383_),
    .A2(_0387_),
    .A3(_0398_),
    .A4(_0400_),
    .B1(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__o22a_1 _2363_ (.A1(\MAC.add.a1[15] ),
    .A2(_0837_),
    .B1(_0380_),
    .B2(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__and3_1 _2364_ (.A(_0482_),
    .B(_0483_),
    .C(_0408_),
    .X(_0411_));
 sky130_fd_sc_hd__or2_1 _2365_ (.A(_0411_),
    .B(_0380_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _2366_ (.A0(\MAC.add.b1[15] ),
    .A1(_0410_),
    .S(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__and3b_1 _2367_ (.A_N(_0809_),
    .B(_0792_),
    .C(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _2368_ (.A(_0414_),
    .X(_0042_));
 sky130_fd_sc_hd__a21o_1 _2369_ (.A1(_0000_),
    .A2(net2),
    .B1(_0002_),
    .X(_0043_));
 sky130_fd_sc_hd__a21o_1 _2370_ (.A1(_0000_),
    .A2(net3),
    .B1(_0009_),
    .X(_0044_));
 sky130_fd_sc_hd__a21o_1 _2371_ (.A1(_0000_),
    .A2(net4),
    .B1(_0010_),
    .X(_0045_));
 sky130_fd_sc_hd__a21o_1 _2372_ (.A1(_0000_),
    .A2(net5),
    .B1(_0011_),
    .X(_0046_));
 sky130_fd_sc_hd__a21o_1 _2373_ (.A1(_0000_),
    .A2(net6),
    .B1(_0012_),
    .X(_0047_));
 sky130_fd_sc_hd__a21o_1 _2374_ (.A1(_0000_),
    .A2(net7),
    .B1(_0013_),
    .X(_0048_));
 sky130_fd_sc_hd__a21o_1 _2375_ (.A1(_0000_),
    .A2(net8),
    .B1(_0014_),
    .X(_0049_));
 sky130_fd_sc_hd__a21o_1 _2376_ (.A1(_0000_),
    .A2(net9),
    .B1(_0015_),
    .X(_0050_));
 sky130_fd_sc_hd__a21o_1 _2377_ (.A1(_0000_),
    .A2(net10),
    .B1(_0016_),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_1 _2378_ (.A1(_0415_),
    .A2(net11),
    .B1(_0017_),
    .X(_0052_));
 sky130_fd_sc_hd__a21o_1 _2379_ (.A1(_0415_),
    .A2(net12),
    .B1(_0003_),
    .X(_0053_));
 sky130_fd_sc_hd__a21o_1 _2380_ (.A1(_0415_),
    .A2(net13),
    .B1(_0004_),
    .X(_0054_));
 sky130_fd_sc_hd__a21o_1 _2381_ (.A1(_0415_),
    .A2(net14),
    .B1(_0005_),
    .X(_0055_));
 sky130_fd_sc_hd__a21o_1 _2382_ (.A1(_0415_),
    .A2(net15),
    .B1(_0006_),
    .X(_0056_));
 sky130_fd_sc_hd__a21o_1 _2383_ (.A1(_0415_),
    .A2(net16),
    .B1(_0007_),
    .X(_0057_));
 sky130_fd_sc_hd__a21o_1 _2384_ (.A1(_0415_),
    .A2(net17),
    .B1(_0008_),
    .X(_0058_));
 sky130_fd_sc_hd__dfrtp_2 _2385_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0018_),
    .RESET_B(net20),
    .Q(\MAC.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2386_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0025_),
    .RESET_B(net20),
    .Q(\MAC.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2387_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0026_),
    .RESET_B(net22),
    .Q(\MAC.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2388_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0027_),
    .RESET_B(net19),
    .Q(\MAC.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2389_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0028_),
    .RESET_B(net19),
    .Q(\MAC.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2390_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0029_),
    .RESET_B(net19),
    .Q(\MAC.b[5] ));
 sky130_fd_sc_hd__dfrtp_4 _2391_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0030_),
    .RESET_B(net22),
    .Q(\MAC.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2392_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0031_),
    .RESET_B(net19),
    .Q(\MAC.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2393_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0032_),
    .RESET_B(net20),
    .Q(\MAC.b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2394_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0033_),
    .RESET_B(net22),
    .Q(\MAC.b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2395_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0019_),
    .RESET_B(net25),
    .Q(\MAC.b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2396_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0020_),
    .RESET_B(net23),
    .Q(\MAC.b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2397_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0021_),
    .RESET_B(net24),
    .Q(\MAC.b[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2398_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0022_),
    .RESET_B(net24),
    .Q(\MAC.b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2399_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0023_),
    .RESET_B(net24),
    .Q(\MAC.b[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2400_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0024_),
    .RESET_B(net22),
    .Q(\MAC.b[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2401_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0002_),
    .RESET_B(net20),
    .Q(\MAC.a[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2402_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0009_),
    .RESET_B(net20),
    .Q(\MAC.a[1] ));
 sky130_fd_sc_hd__dfrtp_4 _2403_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0010_),
    .RESET_B(net22),
    .Q(\MAC.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2404_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0011_),
    .RESET_B(net19),
    .Q(\MAC.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2405_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0012_),
    .RESET_B(net19),
    .Q(\MAC.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2406_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0013_),
    .RESET_B(net19),
    .Q(\MAC.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2407_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0014_),
    .RESET_B(net22),
    .Q(\MAC.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2408_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0015_),
    .RESET_B(net19),
    .Q(\MAC.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2409_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0016_),
    .RESET_B(net20),
    .Q(\MAC.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2410_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0017_),
    .RESET_B(net22),
    .Q(\MAC.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2411_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0003_),
    .RESET_B(net25),
    .Q(\MAC.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2412_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0004_),
    .RESET_B(net24),
    .Q(\MAC.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2413_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0005_),
    .RESET_B(net24),
    .Q(\MAC.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2414_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0006_),
    .RESET_B(net24),
    .Q(\MAC.a[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2415_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0007_),
    .RESET_B(net24),
    .Q(\MAC.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2416_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0008_),
    .RESET_B(net23),
    .Q(\MAC.a[15] ));
 sky130_fd_sc_hd__dfrtp_4 _2417_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0042_),
    .RESET_B(net27),
    .Q(\MAC.add.b1[15] ));
 sky130_fd_sc_hd__dfrtp_4 _2418_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0001_),
    .RESET_B(net28),
    .Q(\wrap2.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2419_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0034_),
    .RESET_B(net28),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfrtp_4 _2420_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0035_),
    .RESET_B(net29),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfrtp_4 _2421_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0036_),
    .RESET_B(net28),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfrtp_4 _2422_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0037_),
    .RESET_B(net28),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__dfrtp_4 _2423_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0038_),
    .RESET_B(net26),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfrtp_4 _2424_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0039_),
    .RESET_B(net26),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfrtp_4 _2425_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0040_),
    .RESET_B(net26),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfrtp_4 _2426_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0041_),
    .RESET_B(net27),
    .Q(uo_out[7]));
 sky130_fd_sc_hd__dfrtp_2 _2427_ (.CLK(clknet_3_6__leaf_clk),
    .D(\MAC.add.c_add[0] ),
    .RESET_B(net27),
    .Q(\MAC.add.b1[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2428_ (.CLK(clknet_3_6__leaf_clk),
    .D(\MAC.add.c_add[1] ),
    .RESET_B(net28),
    .Q(\MAC.add.b1[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2429_ (.CLK(clknet_3_6__leaf_clk),
    .D(\MAC.add.c_add[2] ),
    .RESET_B(net27),
    .Q(\MAC.add.b1[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2430_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.add.c_add[3] ),
    .RESET_B(net27),
    .Q(\MAC.add.b1[3] ));
 sky130_fd_sc_hd__dfrtp_4 _2431_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.add.c_add[4] ),
    .RESET_B(net27),
    .Q(\MAC.add.b1[4] ));
 sky130_fd_sc_hd__dfrtp_2 _2432_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.add.c_add[5] ),
    .RESET_B(net27),
    .Q(\MAC.add.b1[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2433_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.add.c_add[6] ),
    .RESET_B(net27),
    .Q(\MAC.add.b1[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2434_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.add.c_add[7] ),
    .RESET_B(net27),
    .Q(\MAC.add.b1[7] ));
 sky130_fd_sc_hd__dfrtp_4 _2435_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.add.c_add[8] ),
    .RESET_B(net28),
    .Q(\MAC.add.b1[8] ));
 sky130_fd_sc_hd__dfrtp_2 _2436_ (.CLK(clknet_3_6__leaf_clk),
    .D(\MAC.add.c_add[9] ),
    .RESET_B(net28),
    .Q(\MAC.add.b1[9] ));
 sky130_fd_sc_hd__dfrtp_4 _2437_ (.CLK(clknet_3_6__leaf_clk),
    .D(\MAC.add.c_add[10] ),
    .RESET_B(net27),
    .Q(\MAC.add.b1[10] ));
 sky130_fd_sc_hd__dfrtp_4 _2438_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.add.c_add[11] ),
    .RESET_B(net26),
    .Q(\MAC.add.b1[11] ));
 sky130_fd_sc_hd__dfrtp_4 _2439_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.add.c_add[12] ),
    .RESET_B(net26),
    .Q(\MAC.add.b1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2440_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.add.c_add[13] ),
    .RESET_B(net26),
    .Q(\MAC.add.b1[13] ));
 sky130_fd_sc_hd__dfrtp_4 _2441_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.add.c_add[14] ),
    .RESET_B(net26),
    .Q(\MAC.add.b1[14] ));
 sky130_fd_sc_hd__dfrtp_2 _2442_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0000_),
    .RESET_B(net23),
    .Q(\wrap.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2443_ (.CLK(clknet_3_6__leaf_clk),
    .D(\MAC.mul.c_mul1[0] ),
    .RESET_B(net29),
    .Q(\MAC.add.a1[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2444_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[1] ),
    .RESET_B(net21),
    .Q(\MAC.add.a1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2445_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[2] ),
    .RESET_B(net21),
    .Q(\MAC.add.a1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2446_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[3] ),
    .RESET_B(net21),
    .Q(\MAC.add.a1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2447_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[4] ),
    .RESET_B(net21),
    .Q(\MAC.add.a1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2448_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[5] ),
    .RESET_B(net21),
    .Q(\MAC.add.a1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2449_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[6] ),
    .RESET_B(net21),
    .Q(\MAC.add.a1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2450_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[7] ),
    .RESET_B(net21),
    .Q(\MAC.add.a1[7] ));
 sky130_fd_sc_hd__dfrtp_4 _2451_ (.CLK(clknet_3_2__leaf_clk),
    .D(\MAC.mul.c_mul1[8] ),
    .RESET_B(net21),
    .Q(\MAC.add.a1[8] ));
 sky130_fd_sc_hd__dfrtp_2 _2452_ (.CLK(clknet_3_6__leaf_clk),
    .D(\MAC.mul.c_mul1[9] ),
    .RESET_B(net29),
    .Q(\MAC.add.a1[9] ));
 sky130_fd_sc_hd__dfrtp_2 _2453_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.mul.c_mul1[10] ),
    .RESET_B(net29),
    .Q(\MAC.add.a1[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2454_ (.CLK(clknet_3_5__leaf_clk),
    .D(\MAC.mul.c_mul1[11] ),
    .RESET_B(net26),
    .Q(\MAC.add.a1[11] ));
 sky130_fd_sc_hd__dfrtp_4 _2455_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.mul.c_mul1[12] ),
    .RESET_B(net26),
    .Q(\MAC.add.a1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2456_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.mul.c_mul1[13] ),
    .RESET_B(net26),
    .Q(\MAC.add.a1[13] ));
 sky130_fd_sc_hd__dfrtp_2 _2457_ (.CLK(clknet_3_7__leaf_clk),
    .D(\MAC.mul.c_mul1[14] ),
    .RESET_B(net29),
    .Q(\MAC.add.a1[14] ));
 sky130_fd_sc_hd__dfrtp_4 _2458_ (.CLK(clknet_3_6__leaf_clk),
    .D(\MAC.mul.c_mul1[15] ),
    .RESET_B(net29),
    .Q(\MAC.add.a1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2459_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0043_),
    .RESET_B(net22),
    .Q(\wrap.temp_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2460_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0044_),
    .RESET_B(net20),
    .Q(\wrap.temp_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2461_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0045_),
    .RESET_B(net22),
    .Q(\wrap.temp_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2462_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0046_),
    .RESET_B(net20),
    .Q(\wrap.temp_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2463_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0047_),
    .RESET_B(net19),
    .Q(\wrap.temp_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2464_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0048_),
    .RESET_B(net19),
    .Q(\wrap.temp_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2465_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0049_),
    .RESET_B(net22),
    .Q(\wrap.temp_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2466_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0050_),
    .RESET_B(net20),
    .Q(\wrap.temp_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2467_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0051_),
    .RESET_B(net21),
    .Q(\wrap.temp_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2468_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0052_),
    .RESET_B(net23),
    .Q(\wrap.temp_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2469_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0053_),
    .RESET_B(net23),
    .Q(\wrap.temp_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2470_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0054_),
    .RESET_B(net23),
    .Q(\wrap.temp_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2471_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0055_),
    .RESET_B(net23),
    .Q(\wrap.temp_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2472_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0056_),
    .RESET_B(net23),
    .Q(\wrap.temp_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2473_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0057_),
    .RESET_B(net23),
    .Q(\wrap.temp_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2474_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0058_),
    .RESET_B(net23),
    .Q(\wrap.temp_data[15] ));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_45 (.LO(net45));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_542 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(uio_in[2]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(uio_in[3]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(uio_in[4]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(uio_in[5]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(uio_in[6]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(uio_in[7]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 wire18 (.A(_0504_),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(net1),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 fanout22 (.A(net25),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(net25),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 fanout25 (.A(net1),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 fanout26 (.A(net29),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(net1),
    .X(net29));
 sky130_fd_sc_hd__conb_1 tt_um_dlfloatmac_30 (.LO(net30));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload2 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload3 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload4 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload5 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload6 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\wrap.temp_data[0] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\wrap2.state[0] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\wrap.temp_data[10] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\wrap.temp_data[15] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\wrap.temp_data[2] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\wrap.temp_data[9] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\wrap.temp_data[8] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\wrap.temp_data[6] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\wrap.temp_data[1] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\wrap.temp_data[7] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\wrap.temp_data[5] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\wrap.temp_data[11] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\wrap.temp_data[12] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\wrap.temp_data[13] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\wrap.temp_data[4] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\wrap.temp_data[3] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\wrap.temp_data[14] ),
    .X(net62));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_331 ();
 assign uio_oe[0] = net30;
 assign uio_oe[1] = net31;
 assign uio_oe[2] = net32;
 assign uio_oe[3] = net33;
 assign uio_oe[4] = net34;
 assign uio_oe[5] = net35;
 assign uio_oe[6] = net36;
 assign uio_oe[7] = net37;
 assign uio_out[0] = net38;
 assign uio_out[1] = net39;
 assign uio_out[2] = net40;
 assign uio_out[3] = net41;
 assign uio_out[4] = net42;
 assign uio_out[5] = net43;
 assign uio_out[6] = net44;
 assign uio_out[7] = net45;
endmodule
